magic
tech scmos
timestamp 1638537824
<< nwell >>
rect 2 -2 81 27
<< ntransistor >>
rect 13 -45 15 -41
rect 29 -45 31 -41
rect 49 -45 51 -41
rect 68 -45 70 -41
<< ptransistor >>
rect 13 4 15 17
rect 29 4 31 17
rect 49 4 51 17
rect 68 4 70 17
<< ndiffusion >>
rect 12 -45 13 -41
rect 15 -45 16 -41
rect 28 -45 29 -41
rect 31 -45 32 -41
rect 48 -45 49 -41
rect 51 -45 52 -41
rect 67 -45 68 -41
rect 70 -45 71 -41
<< pdiffusion >>
rect 12 4 13 17
rect 15 4 16 17
rect 28 4 29 17
rect 31 4 32 17
rect 48 4 49 17
rect 51 4 52 17
rect 67 4 68 17
rect 70 4 71 17
<< ndcontact >>
rect 8 -45 12 -41
rect 16 -45 20 -41
rect 24 -45 28 -41
rect 32 -45 36 -41
rect 44 -45 48 -41
rect 52 -45 56 -41
rect 63 -45 67 -41
rect 71 -45 75 -41
<< pdcontact >>
rect 8 4 12 17
rect 16 4 20 17
rect 24 4 28 17
rect 32 4 36 17
rect 44 4 48 17
rect 52 4 56 17
rect 63 4 67 17
rect 71 4 75 17
<< polysilicon >>
rect 13 17 15 21
rect 29 17 31 21
rect 49 17 51 21
rect 68 17 70 20
rect 13 -41 15 4
rect 29 -41 31 4
rect 49 -41 51 4
rect 68 -41 70 4
rect 13 -49 15 -45
rect 29 -49 31 -45
rect 49 -50 51 -45
rect 68 -48 70 -45
<< polycontact >>
rect 8 -33 13 -28
rect 24 -8 29 -4
rect 45 -28 49 -23
rect 64 -38 68 -33
<< metal1 >>
rect 2 26 81 30
rect 8 17 12 26
rect 24 17 28 26
rect 44 20 83 23
rect 44 17 48 20
rect 63 17 67 20
rect 3 -28 8 -23
rect 16 -33 20 4
rect 24 -18 29 -13
rect 32 -33 36 4
rect 52 -8 56 4
rect 71 -8 75 4
rect 52 -16 56 -13
rect 52 -20 75 -16
rect 52 -33 56 -29
rect 32 -37 56 -33
rect 16 -41 20 -38
rect 32 -41 36 -37
rect 52 -41 56 -37
rect 71 -41 75 -20
rect 79 -21 83 20
rect 79 -26 85 -21
rect 8 -54 12 -45
rect 24 -54 28 -45
rect 44 -48 48 -45
rect 63 -48 67 -45
rect 79 -48 83 -26
rect 44 -51 83 -48
rect -1 -58 81 -54
<< m2contact >>
rect 8 -28 13 -23
rect 24 -13 29 -8
rect 52 -13 57 -8
rect 71 -13 76 -8
rect 40 -28 45 -23
rect 52 -29 57 -24
rect 16 -38 21 -33
rect 59 -38 64 -33
<< metal2 >>
rect 29 -13 52 -8
rect 63 -13 71 -8
rect 63 -14 76 -13
rect 63 -18 67 -14
rect 52 -22 67 -18
rect 13 -28 40 -23
rect 52 -24 57 -22
rect 21 -38 59 -33
<< labels >>
rlabel metal1 80 -26 85 -21 7 out
rlabel metal1 24 -18 29 -13 1 b
rlabel metal1 3 -28 8 -23 1 a
rlabel metal1 22 28 29 29 5 vdd
rlabel metal1 29 -57 36 -56 1 gnd
<< end >>
