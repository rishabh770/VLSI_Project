magic
tech scmos
timestamp 1638792615
<< nwell >>
rect 19 -23 154 1
rect 211 0 352 1
rect 211 -23 394 0
rect 19 -94 154 -70
rect 209 -71 451 -70
rect 504 -71 540 -70
rect 209 -94 494 -71
rect 500 -94 582 -71
rect 19 -165 154 -141
rect 221 -142 539 -141
rect 221 -165 581 -142
rect 18 -236 153 -212
rect 221 -236 618 -212
<< ntransistor >>
rect 30 -56 32 -52
rect 46 -56 48 -52
rect 62 -56 64 -52
rect 83 -56 85 -52
rect 102 -56 104 -52
rect 122 -56 124 -52
rect 141 -56 143 -52
rect 223 -56 225 -52
rect 239 -56 241 -52
rect 255 -56 257 -52
rect 271 -56 273 -52
rect 291 -56 293 -52
rect 307 -56 309 -52
rect 323 -56 325 -52
rect 341 -56 343 -52
rect 360 -56 362 -52
rect 380 -56 382 -52
rect 30 -127 32 -123
rect 46 -127 48 -123
rect 62 -127 64 -123
rect 83 -127 85 -123
rect 102 -127 104 -123
rect 122 -127 124 -123
rect 141 -127 143 -123
rect 221 -127 223 -123
rect 241 -127 243 -123
rect 257 -127 259 -123
rect 273 -127 275 -123
rect 289 -127 291 -123
rect 305 -127 307 -123
rect 321 -127 323 -123
rect 340 -127 342 -123
rect 359 -127 361 -123
rect 375 -127 377 -123
rect 391 -127 393 -123
rect 407 -127 409 -123
rect 423 -127 425 -123
rect 441 -127 443 -123
rect 460 -127 462 -123
rect 480 -127 482 -123
rect 511 -127 513 -123
rect 529 -127 531 -123
rect 548 -127 550 -123
rect 568 -127 570 -123
rect 30 -198 32 -194
rect 46 -198 48 -194
rect 62 -198 64 -194
rect 83 -198 85 -194
rect 102 -198 104 -194
rect 122 -198 124 -194
rect 141 -198 143 -194
rect 232 -198 234 -194
rect 248 -198 250 -194
rect 264 -198 266 -194
rect 280 -198 282 -194
rect 296 -198 298 -194
rect 315 -198 317 -194
rect 331 -198 333 -194
rect 347 -198 349 -194
rect 363 -198 365 -194
rect 382 -198 384 -194
rect 398 -198 400 -194
rect 414 -198 416 -194
rect 430 -198 432 -194
rect 446 -198 448 -194
rect 462 -198 464 -194
rect 478 -198 480 -194
rect 494 -198 496 -194
rect 510 -198 512 -194
rect 528 -198 530 -194
rect 547 -198 549 -194
rect 567 -198 569 -194
rect 29 -269 31 -265
rect 45 -269 47 -265
rect 61 -269 63 -265
rect 82 -269 84 -265
rect 101 -269 103 -265
rect 121 -269 123 -265
rect 140 -269 142 -265
rect 232 -269 234 -265
rect 248 -269 250 -265
rect 264 -269 266 -265
rect 280 -269 282 -265
rect 296 -269 298 -265
rect 312 -269 314 -265
rect 328 -269 330 -265
rect 344 -269 346 -265
rect 360 -269 362 -265
rect 376 -269 378 -265
rect 392 -269 394 -265
rect 412 -269 414 -265
rect 428 -269 430 -265
rect 444 -269 446 -265
rect 460 -269 462 -265
rect 477 -269 479 -265
rect 493 -269 495 -265
rect 509 -269 511 -265
rect 525 -269 527 -265
rect 541 -269 543 -265
rect 557 -269 559 -265
rect 573 -269 575 -265
rect 589 -269 591 -265
rect 605 -269 607 -265
<< ptransistor >>
rect 30 -16 32 -7
rect 46 -16 48 -7
rect 62 -16 64 -7
rect 83 -16 85 -7
rect 102 -16 104 -7
rect 122 -16 124 -7
rect 141 -16 143 -7
rect 223 -16 225 -7
rect 239 -16 241 -7
rect 255 -16 257 -7
rect 271 -16 273 -7
rect 291 -16 293 -7
rect 307 -16 309 -7
rect 323 -16 325 -7
rect 341 -16 343 -7
rect 360 -16 362 -7
rect 380 -16 382 -7
rect 30 -87 32 -78
rect 46 -87 48 -78
rect 62 -87 64 -78
rect 83 -87 85 -78
rect 102 -87 104 -78
rect 122 -87 124 -78
rect 141 -87 143 -78
rect 221 -87 223 -78
rect 241 -87 243 -78
rect 257 -87 259 -78
rect 273 -87 275 -78
rect 289 -87 291 -78
rect 305 -87 307 -78
rect 321 -87 323 -78
rect 340 -87 342 -78
rect 359 -87 361 -78
rect 375 -87 377 -78
rect 391 -87 393 -78
rect 407 -87 409 -78
rect 423 -87 425 -78
rect 441 -87 443 -78
rect 460 -87 462 -78
rect 480 -87 482 -78
rect 511 -87 513 -78
rect 529 -87 531 -78
rect 548 -87 550 -78
rect 568 -87 570 -78
rect 30 -158 32 -149
rect 46 -158 48 -149
rect 62 -158 64 -149
rect 83 -158 85 -149
rect 102 -158 104 -149
rect 122 -158 124 -149
rect 141 -158 143 -149
rect 232 -158 234 -149
rect 248 -158 250 -149
rect 264 -158 266 -149
rect 280 -158 282 -149
rect 296 -158 298 -149
rect 315 -158 317 -149
rect 331 -158 333 -149
rect 347 -158 349 -149
rect 363 -158 365 -149
rect 382 -158 384 -149
rect 398 -158 400 -149
rect 414 -158 416 -149
rect 430 -158 432 -149
rect 446 -158 448 -149
rect 462 -158 464 -149
rect 478 -158 480 -149
rect 494 -158 496 -149
rect 510 -158 512 -149
rect 528 -158 530 -149
rect 547 -158 549 -149
rect 567 -158 569 -149
rect 29 -229 31 -220
rect 45 -229 47 -220
rect 61 -229 63 -220
rect 82 -229 84 -220
rect 101 -229 103 -220
rect 121 -229 123 -220
rect 140 -229 142 -220
rect 232 -229 234 -220
rect 248 -229 250 -220
rect 264 -229 266 -220
rect 280 -229 282 -220
rect 296 -229 298 -220
rect 312 -229 314 -220
rect 328 -229 330 -220
rect 344 -229 346 -220
rect 360 -229 362 -220
rect 376 -229 378 -220
rect 392 -229 394 -220
rect 412 -229 414 -220
rect 428 -229 430 -220
rect 444 -229 446 -220
rect 460 -229 462 -220
rect 477 -229 479 -220
rect 493 -229 495 -220
rect 509 -229 511 -220
rect 525 -229 527 -220
rect 541 -229 543 -220
rect 557 -229 559 -220
rect 573 -229 575 -220
rect 589 -229 591 -220
rect 605 -229 607 -220
<< ndiffusion >>
rect 29 -56 30 -52
rect 32 -56 33 -52
rect 45 -56 46 -52
rect 48 -56 49 -52
rect 61 -56 62 -52
rect 64 -56 65 -52
rect 82 -56 83 -52
rect 85 -56 86 -52
rect 101 -56 102 -52
rect 104 -56 105 -52
rect 121 -56 122 -52
rect 124 -56 125 -52
rect 140 -56 141 -52
rect 143 -56 144 -52
rect 222 -56 223 -52
rect 225 -56 226 -52
rect 238 -56 239 -52
rect 241 -56 242 -52
rect 254 -56 255 -52
rect 257 -56 258 -52
rect 270 -56 271 -52
rect 273 -56 274 -52
rect 290 -56 291 -52
rect 293 -56 294 -52
rect 306 -56 307 -52
rect 309 -56 310 -52
rect 322 -56 323 -52
rect 325 -56 326 -52
rect 340 -56 341 -52
rect 343 -56 344 -52
rect 359 -56 360 -52
rect 362 -56 363 -52
rect 379 -56 380 -52
rect 382 -56 383 -52
rect 29 -127 30 -123
rect 32 -127 33 -123
rect 45 -127 46 -123
rect 48 -127 49 -123
rect 61 -127 62 -123
rect 64 -127 65 -123
rect 82 -127 83 -123
rect 85 -127 86 -123
rect 101 -127 102 -123
rect 104 -127 105 -123
rect 121 -127 122 -123
rect 124 -127 125 -123
rect 140 -127 141 -123
rect 143 -127 144 -123
rect 220 -127 221 -123
rect 223 -127 224 -123
rect 240 -127 241 -123
rect 243 -127 244 -123
rect 256 -127 257 -123
rect 259 -127 260 -123
rect 272 -127 273 -123
rect 275 -127 276 -123
rect 288 -127 289 -123
rect 291 -127 292 -123
rect 304 -127 305 -123
rect 307 -127 308 -123
rect 320 -127 321 -123
rect 323 -127 324 -123
rect 339 -127 340 -123
rect 342 -127 343 -123
rect 358 -127 359 -123
rect 361 -127 362 -123
rect 374 -127 375 -123
rect 377 -127 378 -123
rect 390 -127 391 -123
rect 393 -127 394 -123
rect 406 -127 407 -123
rect 409 -127 410 -123
rect 422 -127 423 -123
rect 425 -127 426 -123
rect 440 -127 441 -123
rect 443 -127 444 -123
rect 459 -127 460 -123
rect 462 -127 463 -123
rect 479 -127 480 -123
rect 482 -127 483 -123
rect 510 -127 511 -123
rect 513 -127 514 -123
rect 528 -127 529 -123
rect 531 -127 532 -123
rect 547 -127 548 -123
rect 550 -127 551 -123
rect 567 -127 568 -123
rect 570 -127 571 -123
rect 29 -198 30 -194
rect 32 -198 33 -194
rect 45 -198 46 -194
rect 48 -198 49 -194
rect 61 -198 62 -194
rect 64 -198 65 -194
rect 82 -198 83 -194
rect 85 -198 86 -194
rect 101 -198 102 -194
rect 104 -198 105 -194
rect 121 -198 122 -194
rect 124 -198 125 -194
rect 140 -198 141 -194
rect 143 -198 144 -194
rect 231 -198 232 -194
rect 234 -198 235 -194
rect 247 -198 248 -194
rect 250 -198 251 -194
rect 263 -198 264 -194
rect 266 -198 267 -194
rect 279 -198 280 -194
rect 282 -198 283 -194
rect 295 -198 296 -194
rect 298 -198 299 -194
rect 314 -198 315 -194
rect 317 -198 318 -194
rect 330 -198 331 -194
rect 333 -198 334 -194
rect 346 -198 347 -194
rect 349 -198 350 -194
rect 362 -198 363 -194
rect 365 -198 366 -194
rect 381 -198 382 -194
rect 384 -198 385 -194
rect 397 -198 398 -194
rect 400 -198 401 -194
rect 413 -198 414 -194
rect 416 -198 417 -194
rect 429 -198 430 -194
rect 432 -198 433 -194
rect 445 -198 446 -194
rect 448 -198 449 -194
rect 461 -198 462 -194
rect 464 -198 465 -194
rect 477 -198 478 -194
rect 480 -198 481 -194
rect 493 -198 494 -194
rect 496 -198 497 -194
rect 509 -198 510 -194
rect 512 -198 513 -194
rect 527 -198 528 -194
rect 530 -198 531 -194
rect 546 -198 547 -194
rect 549 -198 550 -194
rect 566 -198 567 -194
rect 569 -198 570 -194
rect 28 -269 29 -265
rect 31 -269 32 -265
rect 44 -269 45 -265
rect 47 -269 48 -265
rect 60 -269 61 -265
rect 63 -269 64 -265
rect 81 -269 82 -265
rect 84 -269 85 -265
rect 100 -269 101 -265
rect 103 -269 104 -265
rect 120 -269 121 -265
rect 123 -269 124 -265
rect 139 -269 140 -265
rect 142 -269 143 -265
rect 231 -269 232 -265
rect 234 -269 235 -265
rect 247 -269 248 -265
rect 250 -269 251 -265
rect 263 -269 264 -265
rect 266 -269 267 -265
rect 279 -269 280 -265
rect 282 -269 283 -265
rect 295 -269 296 -265
rect 298 -269 299 -265
rect 311 -269 312 -265
rect 314 -269 315 -265
rect 327 -269 328 -265
rect 330 -269 331 -265
rect 343 -269 344 -265
rect 346 -269 347 -265
rect 359 -269 360 -265
rect 362 -269 363 -265
rect 375 -269 376 -265
rect 378 -269 379 -265
rect 391 -269 392 -265
rect 394 -269 395 -265
rect 411 -269 412 -265
rect 414 -269 415 -265
rect 427 -269 428 -265
rect 430 -269 431 -265
rect 443 -269 444 -265
rect 446 -269 447 -265
rect 459 -269 460 -265
rect 462 -269 463 -265
rect 476 -269 477 -265
rect 479 -269 480 -265
rect 492 -269 493 -265
rect 495 -269 496 -265
rect 508 -269 509 -265
rect 511 -269 512 -265
rect 524 -269 525 -265
rect 527 -269 528 -265
rect 540 -269 541 -265
rect 543 -269 544 -265
rect 556 -269 557 -265
rect 559 -269 560 -265
rect 572 -269 573 -265
rect 575 -269 576 -265
rect 588 -269 589 -265
rect 591 -269 592 -265
rect 604 -269 605 -265
rect 607 -269 608 -265
<< pdiffusion >>
rect 29 -16 30 -7
rect 32 -16 33 -7
rect 45 -16 46 -7
rect 48 -16 49 -7
rect 61 -16 62 -7
rect 64 -16 65 -7
rect 82 -16 83 -7
rect 85 -16 86 -7
rect 101 -16 102 -7
rect 104 -16 105 -7
rect 121 -16 122 -7
rect 124 -16 125 -7
rect 140 -16 141 -7
rect 143 -16 144 -7
rect 222 -16 223 -7
rect 225 -16 226 -7
rect 238 -16 239 -7
rect 241 -16 242 -7
rect 254 -16 255 -7
rect 257 -16 258 -7
rect 270 -16 271 -7
rect 273 -16 274 -7
rect 290 -16 291 -7
rect 293 -16 294 -7
rect 306 -16 307 -7
rect 309 -16 310 -7
rect 322 -16 323 -7
rect 325 -16 326 -7
rect 340 -16 341 -7
rect 343 -16 344 -7
rect 359 -16 360 -7
rect 362 -16 363 -7
rect 379 -16 380 -7
rect 382 -16 383 -7
rect 29 -87 30 -78
rect 32 -87 33 -78
rect 45 -87 46 -78
rect 48 -87 49 -78
rect 61 -87 62 -78
rect 64 -87 65 -78
rect 82 -87 83 -78
rect 85 -87 86 -78
rect 101 -87 102 -78
rect 104 -87 105 -78
rect 121 -87 122 -78
rect 124 -87 125 -78
rect 140 -87 141 -78
rect 143 -87 144 -78
rect 220 -87 221 -78
rect 223 -87 224 -78
rect 240 -87 241 -78
rect 243 -87 244 -78
rect 256 -87 257 -78
rect 259 -87 260 -78
rect 272 -87 273 -78
rect 275 -87 276 -78
rect 288 -87 289 -78
rect 291 -87 292 -78
rect 304 -87 305 -78
rect 307 -87 308 -78
rect 320 -87 321 -78
rect 323 -87 324 -78
rect 339 -87 340 -78
rect 342 -87 343 -78
rect 358 -87 359 -78
rect 361 -87 362 -78
rect 374 -87 375 -78
rect 377 -87 378 -78
rect 390 -87 391 -78
rect 393 -87 394 -78
rect 406 -87 407 -78
rect 409 -87 410 -78
rect 422 -87 423 -78
rect 425 -87 426 -78
rect 440 -87 441 -78
rect 443 -87 444 -78
rect 459 -87 460 -78
rect 462 -87 463 -78
rect 479 -87 480 -78
rect 482 -87 483 -78
rect 510 -87 511 -78
rect 513 -87 514 -78
rect 528 -87 529 -78
rect 531 -87 532 -78
rect 547 -87 548 -78
rect 550 -87 551 -78
rect 567 -87 568 -78
rect 570 -87 571 -78
rect 29 -158 30 -149
rect 32 -158 33 -149
rect 45 -158 46 -149
rect 48 -158 49 -149
rect 61 -158 62 -149
rect 64 -158 65 -149
rect 82 -158 83 -149
rect 85 -158 86 -149
rect 101 -158 102 -149
rect 104 -158 105 -149
rect 121 -158 122 -149
rect 124 -158 125 -149
rect 140 -158 141 -149
rect 143 -158 144 -149
rect 231 -158 232 -149
rect 234 -158 235 -149
rect 247 -158 248 -149
rect 250 -158 251 -149
rect 263 -158 264 -149
rect 266 -158 267 -149
rect 279 -158 280 -149
rect 282 -158 283 -149
rect 295 -158 296 -149
rect 298 -158 299 -149
rect 314 -158 315 -149
rect 317 -158 318 -149
rect 330 -158 331 -149
rect 333 -158 334 -149
rect 346 -158 347 -149
rect 349 -158 350 -149
rect 362 -158 363 -149
rect 365 -158 366 -149
rect 381 -158 382 -149
rect 384 -158 385 -149
rect 397 -158 398 -149
rect 400 -158 401 -149
rect 413 -158 414 -149
rect 416 -158 417 -149
rect 429 -158 430 -149
rect 432 -158 433 -149
rect 445 -158 446 -149
rect 448 -158 449 -149
rect 461 -158 462 -149
rect 464 -158 465 -149
rect 477 -158 478 -149
rect 480 -158 481 -149
rect 493 -158 494 -149
rect 496 -158 497 -149
rect 509 -158 510 -149
rect 512 -158 513 -149
rect 527 -158 528 -149
rect 530 -158 531 -149
rect 546 -158 547 -149
rect 549 -158 550 -149
rect 566 -158 567 -149
rect 569 -158 570 -149
rect 28 -229 29 -220
rect 31 -229 32 -220
rect 44 -229 45 -220
rect 47 -229 48 -220
rect 60 -229 61 -220
rect 63 -229 64 -220
rect 81 -229 82 -220
rect 84 -229 85 -220
rect 100 -229 101 -220
rect 103 -229 104 -220
rect 120 -229 121 -220
rect 123 -229 124 -220
rect 139 -229 140 -220
rect 142 -229 143 -220
rect 231 -229 232 -220
rect 234 -229 235 -220
rect 247 -229 248 -220
rect 250 -229 251 -220
rect 263 -229 264 -220
rect 266 -229 267 -220
rect 279 -229 280 -220
rect 282 -229 283 -220
rect 295 -229 296 -220
rect 298 -229 299 -220
rect 311 -229 312 -220
rect 314 -229 315 -220
rect 327 -229 328 -220
rect 330 -229 331 -220
rect 343 -229 344 -220
rect 346 -229 347 -220
rect 359 -229 360 -220
rect 362 -229 363 -220
rect 375 -229 376 -220
rect 378 -229 379 -220
rect 391 -229 392 -220
rect 394 -229 395 -220
rect 411 -229 412 -220
rect 414 -229 415 -220
rect 427 -229 428 -220
rect 430 -229 431 -220
rect 443 -229 444 -220
rect 446 -229 447 -220
rect 459 -229 460 -220
rect 462 -229 463 -220
rect 476 -229 477 -220
rect 479 -229 480 -220
rect 492 -229 493 -220
rect 495 -229 496 -220
rect 508 -229 509 -220
rect 511 -229 512 -220
rect 524 -229 525 -220
rect 527 -229 528 -220
rect 540 -229 541 -220
rect 543 -229 544 -220
rect 556 -229 557 -220
rect 559 -229 560 -220
rect 572 -229 573 -220
rect 575 -229 576 -220
rect 588 -229 589 -220
rect 591 -229 592 -220
rect 604 -229 605 -220
rect 607 -229 608 -220
<< ndcontact >>
rect 25 -56 29 -52
rect 33 -56 37 -52
rect 41 -56 45 -52
rect 49 -56 53 -52
rect 57 -56 61 -52
rect 65 -56 69 -52
rect 78 -56 82 -52
rect 86 -56 90 -52
rect 97 -56 101 -52
rect 105 -56 109 -52
rect 117 -56 121 -52
rect 125 -56 129 -52
rect 136 -56 140 -52
rect 144 -56 148 -52
rect 218 -56 222 -52
rect 226 -56 230 -52
rect 234 -56 238 -52
rect 242 -56 246 -52
rect 250 -56 254 -52
rect 258 -56 262 -52
rect 266 -56 270 -52
rect 274 -56 278 -52
rect 286 -56 290 -52
rect 294 -56 298 -52
rect 302 -56 306 -52
rect 310 -56 314 -52
rect 318 -56 322 -52
rect 326 -56 330 -52
rect 336 -56 340 -52
rect 344 -56 348 -52
rect 355 -56 359 -52
rect 363 -56 367 -52
rect 375 -56 379 -52
rect 383 -56 387 -52
rect 25 -127 29 -123
rect 33 -127 37 -123
rect 41 -127 45 -123
rect 49 -127 53 -123
rect 57 -127 61 -123
rect 65 -127 69 -123
rect 78 -127 82 -123
rect 86 -127 90 -123
rect 97 -127 101 -123
rect 105 -127 109 -123
rect 117 -127 121 -123
rect 125 -127 129 -123
rect 136 -127 140 -123
rect 144 -127 148 -123
rect 216 -127 220 -123
rect 224 -127 228 -123
rect 236 -127 240 -123
rect 244 -127 248 -123
rect 252 -127 256 -123
rect 260 -127 264 -123
rect 268 -127 272 -123
rect 276 -127 280 -123
rect 284 -127 288 -123
rect 292 -127 296 -123
rect 300 -127 304 -123
rect 308 -127 312 -123
rect 316 -127 320 -123
rect 324 -127 328 -123
rect 335 -127 339 -123
rect 343 -127 347 -123
rect 354 -127 358 -123
rect 362 -127 366 -123
rect 370 -127 374 -123
rect 378 -127 382 -123
rect 386 -127 390 -123
rect 394 -127 398 -123
rect 402 -127 406 -123
rect 410 -127 414 -123
rect 418 -127 422 -123
rect 426 -127 430 -123
rect 436 -127 440 -123
rect 444 -127 448 -123
rect 455 -127 459 -123
rect 463 -127 467 -123
rect 475 -127 479 -123
rect 483 -127 487 -123
rect 506 -127 510 -123
rect 514 -127 518 -123
rect 524 -127 528 -123
rect 532 -127 536 -123
rect 543 -127 547 -123
rect 551 -127 555 -123
rect 563 -127 567 -123
rect 571 -127 575 -123
rect 25 -198 29 -194
rect 33 -198 37 -194
rect 41 -198 45 -194
rect 49 -198 53 -194
rect 57 -198 61 -194
rect 65 -198 69 -194
rect 78 -198 82 -194
rect 86 -198 90 -194
rect 97 -198 101 -194
rect 105 -198 109 -194
rect 117 -198 121 -194
rect 125 -198 129 -194
rect 136 -198 140 -194
rect 144 -198 148 -194
rect 227 -198 231 -194
rect 235 -198 239 -194
rect 243 -198 247 -194
rect 251 -198 255 -194
rect 259 -198 263 -194
rect 267 -198 271 -194
rect 275 -198 279 -194
rect 283 -198 287 -194
rect 291 -198 295 -194
rect 299 -198 303 -194
rect 310 -198 314 -194
rect 318 -198 322 -194
rect 326 -198 330 -194
rect 334 -198 338 -194
rect 342 -198 346 -194
rect 350 -198 354 -194
rect 358 -198 362 -194
rect 366 -198 370 -194
rect 377 -198 381 -194
rect 385 -198 389 -194
rect 393 -198 397 -194
rect 401 -198 405 -194
rect 409 -198 413 -194
rect 417 -198 421 -194
rect 425 -198 429 -194
rect 433 -198 437 -194
rect 441 -198 445 -194
rect 449 -198 453 -194
rect 457 -198 461 -194
rect 465 -198 469 -194
rect 473 -198 477 -194
rect 481 -198 485 -194
rect 489 -198 493 -194
rect 497 -198 501 -194
rect 505 -198 509 -194
rect 513 -198 517 -194
rect 523 -198 527 -194
rect 531 -198 535 -194
rect 542 -198 546 -194
rect 550 -198 554 -194
rect 562 -198 566 -194
rect 570 -198 574 -194
rect 24 -269 28 -265
rect 32 -269 36 -265
rect 40 -269 44 -265
rect 48 -269 52 -265
rect 56 -269 60 -265
rect 64 -269 68 -265
rect 77 -269 81 -265
rect 85 -269 89 -265
rect 96 -269 100 -265
rect 104 -269 108 -265
rect 116 -269 120 -265
rect 124 -269 128 -265
rect 135 -269 139 -265
rect 143 -269 147 -265
rect 227 -269 231 -265
rect 235 -269 239 -265
rect 243 -269 247 -265
rect 251 -269 255 -265
rect 259 -269 263 -265
rect 267 -269 271 -265
rect 275 -269 279 -265
rect 283 -269 287 -265
rect 291 -269 295 -265
rect 299 -269 303 -265
rect 307 -269 311 -265
rect 315 -269 319 -265
rect 323 -269 327 -265
rect 331 -269 335 -265
rect 339 -269 343 -265
rect 347 -269 351 -265
rect 355 -269 359 -265
rect 363 -269 367 -265
rect 371 -269 375 -265
rect 379 -269 383 -265
rect 387 -269 391 -265
rect 395 -269 399 -265
rect 407 -269 411 -265
rect 415 -269 419 -265
rect 423 -269 427 -265
rect 431 -269 435 -265
rect 439 -269 443 -265
rect 447 -269 451 -265
rect 455 -269 459 -265
rect 463 -269 467 -265
rect 472 -269 476 -265
rect 480 -269 484 -265
rect 488 -269 492 -265
rect 496 -269 500 -265
rect 504 -269 508 -265
rect 512 -269 516 -265
rect 520 -269 524 -265
rect 528 -269 532 -265
rect 536 -269 540 -265
rect 544 -269 548 -265
rect 552 -269 556 -265
rect 560 -269 564 -265
rect 568 -269 572 -265
rect 576 -269 580 -265
rect 584 -269 588 -265
rect 592 -269 596 -265
rect 600 -269 604 -265
rect 608 -269 612 -265
<< pdcontact >>
rect 25 -16 29 -7
rect 33 -16 37 -7
rect 41 -16 45 -7
rect 49 -16 53 -7
rect 57 -16 61 -7
rect 65 -16 69 -7
rect 78 -16 82 -7
rect 86 -16 90 -7
rect 97 -16 101 -7
rect 105 -16 109 -7
rect 117 -16 121 -7
rect 125 -16 129 -7
rect 136 -16 140 -7
rect 144 -16 148 -7
rect 218 -16 222 -7
rect 226 -16 230 -7
rect 234 -16 238 -7
rect 242 -16 246 -7
rect 250 -16 254 -7
rect 258 -16 262 -7
rect 266 -16 270 -7
rect 274 -16 278 -7
rect 286 -16 290 -7
rect 294 -16 298 -7
rect 302 -16 306 -7
rect 310 -16 314 -7
rect 318 -16 322 -7
rect 326 -16 330 -7
rect 336 -16 340 -7
rect 344 -16 348 -7
rect 355 -16 359 -7
rect 363 -16 367 -7
rect 375 -16 379 -7
rect 383 -16 387 -7
rect 25 -87 29 -78
rect 33 -87 37 -78
rect 41 -87 45 -78
rect 49 -87 53 -78
rect 57 -87 61 -78
rect 65 -87 69 -78
rect 78 -87 82 -78
rect 86 -87 90 -78
rect 97 -87 101 -78
rect 105 -87 109 -78
rect 117 -87 121 -78
rect 125 -87 129 -78
rect 136 -87 140 -78
rect 144 -87 148 -78
rect 216 -87 220 -78
rect 224 -87 228 -78
rect 236 -87 240 -78
rect 244 -87 248 -78
rect 252 -87 256 -78
rect 260 -87 264 -78
rect 268 -87 272 -78
rect 276 -87 280 -78
rect 284 -87 288 -78
rect 292 -87 296 -78
rect 300 -87 304 -78
rect 308 -87 312 -78
rect 316 -87 320 -78
rect 324 -87 328 -78
rect 335 -87 339 -78
rect 343 -87 347 -78
rect 354 -87 358 -78
rect 362 -87 366 -78
rect 370 -87 374 -78
rect 378 -87 382 -78
rect 386 -87 390 -78
rect 394 -87 398 -78
rect 402 -87 406 -78
rect 410 -87 414 -78
rect 418 -87 422 -78
rect 426 -87 430 -78
rect 436 -87 440 -78
rect 444 -87 448 -78
rect 455 -87 459 -78
rect 463 -87 467 -78
rect 475 -87 479 -78
rect 483 -87 487 -78
rect 506 -87 510 -78
rect 514 -87 518 -78
rect 524 -87 528 -78
rect 532 -87 536 -78
rect 543 -87 547 -78
rect 551 -87 555 -78
rect 563 -87 567 -78
rect 571 -87 575 -78
rect 25 -158 29 -149
rect 33 -158 37 -149
rect 41 -158 45 -149
rect 49 -158 53 -149
rect 57 -158 61 -149
rect 65 -158 69 -149
rect 78 -158 82 -149
rect 86 -158 90 -149
rect 97 -158 101 -149
rect 105 -158 109 -149
rect 117 -158 121 -149
rect 125 -158 129 -149
rect 136 -158 140 -149
rect 144 -158 148 -149
rect 227 -158 231 -149
rect 235 -158 239 -149
rect 243 -158 247 -149
rect 251 -158 255 -149
rect 259 -158 263 -149
rect 267 -158 271 -149
rect 275 -158 279 -149
rect 283 -158 287 -149
rect 291 -158 295 -149
rect 299 -158 303 -149
rect 310 -158 314 -149
rect 318 -158 322 -149
rect 326 -158 330 -149
rect 334 -158 338 -149
rect 342 -158 346 -149
rect 350 -158 354 -149
rect 358 -158 362 -149
rect 366 -158 370 -149
rect 377 -158 381 -149
rect 385 -158 389 -149
rect 393 -158 397 -149
rect 401 -158 405 -149
rect 409 -158 413 -149
rect 417 -158 421 -149
rect 425 -158 429 -149
rect 433 -158 437 -149
rect 441 -158 445 -149
rect 449 -158 453 -149
rect 457 -158 461 -149
rect 465 -158 469 -149
rect 473 -158 477 -149
rect 481 -158 485 -149
rect 489 -158 493 -149
rect 497 -158 501 -149
rect 505 -158 509 -149
rect 513 -158 517 -149
rect 523 -158 527 -149
rect 531 -158 535 -149
rect 542 -158 546 -149
rect 550 -158 554 -149
rect 562 -158 566 -149
rect 570 -158 574 -149
rect 24 -229 28 -220
rect 32 -229 36 -220
rect 40 -229 44 -220
rect 48 -229 52 -220
rect 56 -229 60 -220
rect 64 -229 68 -220
rect 77 -229 81 -220
rect 85 -229 89 -220
rect 96 -229 100 -220
rect 104 -229 108 -220
rect 116 -229 120 -220
rect 124 -229 128 -220
rect 135 -229 139 -220
rect 143 -229 147 -220
rect 227 -229 231 -220
rect 235 -229 239 -220
rect 243 -229 247 -220
rect 251 -229 255 -220
rect 259 -229 263 -220
rect 267 -229 271 -220
rect 275 -229 279 -220
rect 283 -229 287 -220
rect 291 -229 295 -220
rect 299 -229 303 -220
rect 307 -229 311 -220
rect 315 -229 319 -220
rect 323 -229 327 -220
rect 331 -229 335 -220
rect 339 -229 343 -220
rect 347 -229 351 -220
rect 355 -229 359 -220
rect 363 -229 367 -220
rect 371 -229 375 -220
rect 379 -229 383 -220
rect 387 -229 391 -220
rect 395 -229 399 -220
rect 407 -229 411 -220
rect 415 -229 419 -220
rect 423 -229 427 -220
rect 431 -229 435 -220
rect 439 -229 443 -220
rect 447 -229 451 -220
rect 455 -229 459 -220
rect 463 -229 467 -220
rect 472 -229 476 -220
rect 480 -229 484 -220
rect 488 -229 492 -220
rect 496 -229 500 -220
rect 504 -229 508 -220
rect 512 -229 516 -220
rect 520 -229 524 -220
rect 528 -229 532 -220
rect 536 -229 540 -220
rect 544 -229 548 -220
rect 552 -229 556 -220
rect 560 -229 564 -220
rect 568 -229 572 -220
rect 576 -229 580 -220
rect 584 -229 588 -220
rect 592 -229 596 -220
rect 600 -229 604 -220
rect 608 -229 612 -220
<< polysilicon >>
rect 30 -7 32 -4
rect 46 -7 48 -4
rect 62 -7 64 -4
rect 83 -7 85 -4
rect 102 -7 104 -4
rect 122 -7 124 -4
rect 141 -7 143 -4
rect 223 -7 225 -4
rect 239 -7 241 -4
rect 255 -7 257 -4
rect 271 -7 273 -4
rect 291 -7 293 -4
rect 307 -7 309 -4
rect 323 -7 325 -4
rect 341 -7 343 -4
rect 360 -7 362 -4
rect 380 -7 382 -4
rect 30 -52 32 -16
rect 46 -52 48 -16
rect 62 -52 64 -16
rect 83 -52 85 -16
rect 102 -52 104 -16
rect 122 -52 124 -16
rect 141 -52 143 -16
rect 223 -52 225 -16
rect 239 -52 241 -16
rect 255 -52 257 -16
rect 271 -52 273 -16
rect 291 -52 293 -16
rect 307 -52 309 -16
rect 323 -52 325 -16
rect 341 -52 343 -16
rect 360 -52 362 -16
rect 380 -52 382 -16
rect 30 -59 32 -56
rect 46 -59 48 -56
rect 62 -59 64 -56
rect 83 -59 85 -56
rect 102 -59 104 -56
rect 122 -59 124 -56
rect 141 -59 143 -56
rect 223 -59 225 -56
rect 239 -59 241 -56
rect 255 -59 257 -56
rect 271 -59 273 -56
rect 291 -59 293 -56
rect 307 -59 309 -56
rect 323 -59 325 -56
rect 341 -59 343 -56
rect 360 -59 362 -56
rect 380 -59 382 -56
rect 30 -78 32 -75
rect 46 -78 48 -75
rect 62 -78 64 -75
rect 83 -78 85 -75
rect 102 -78 104 -75
rect 122 -78 124 -75
rect 141 -78 143 -75
rect 221 -78 223 -75
rect 241 -78 243 -75
rect 257 -78 259 -75
rect 273 -78 275 -75
rect 289 -78 291 -75
rect 305 -78 307 -75
rect 321 -78 323 -75
rect 340 -78 342 -75
rect 359 -78 361 -75
rect 375 -78 377 -75
rect 391 -78 393 -75
rect 407 -78 409 -75
rect 423 -78 425 -75
rect 441 -78 443 -75
rect 460 -78 462 -75
rect 480 -78 482 -75
rect 511 -78 513 -75
rect 529 -78 531 -75
rect 548 -78 550 -75
rect 568 -78 570 -75
rect 30 -123 32 -87
rect 46 -123 48 -87
rect 62 -123 64 -87
rect 83 -123 85 -87
rect 102 -123 104 -87
rect 122 -123 124 -87
rect 141 -123 143 -87
rect 221 -123 223 -87
rect 241 -123 243 -87
rect 257 -123 259 -87
rect 273 -123 275 -87
rect 289 -123 291 -87
rect 305 -123 307 -87
rect 321 -123 323 -87
rect 340 -123 342 -87
rect 359 -123 361 -87
rect 375 -123 377 -87
rect 391 -123 393 -87
rect 407 -123 409 -87
rect 423 -123 425 -87
rect 441 -123 443 -87
rect 460 -123 462 -87
rect 480 -123 482 -87
rect 511 -123 513 -87
rect 529 -123 531 -87
rect 548 -123 550 -87
rect 568 -123 570 -87
rect 30 -130 32 -127
rect 46 -130 48 -127
rect 62 -130 64 -127
rect 83 -130 85 -127
rect 102 -130 104 -127
rect 122 -130 124 -127
rect 141 -130 143 -127
rect 221 -130 223 -127
rect 241 -130 243 -127
rect 257 -130 259 -127
rect 273 -130 275 -127
rect 289 -130 291 -127
rect 305 -130 307 -127
rect 321 -130 323 -127
rect 340 -130 342 -127
rect 359 -130 361 -127
rect 375 -130 377 -127
rect 391 -130 393 -127
rect 407 -130 409 -127
rect 423 -130 425 -127
rect 441 -130 443 -127
rect 460 -130 462 -127
rect 480 -130 482 -127
rect 511 -130 513 -127
rect 529 -130 531 -127
rect 548 -130 550 -127
rect 568 -130 570 -127
rect 30 -149 32 -146
rect 46 -149 48 -146
rect 62 -149 64 -146
rect 83 -149 85 -146
rect 102 -149 104 -146
rect 122 -149 124 -146
rect 141 -149 143 -146
rect 232 -149 234 -146
rect 248 -149 250 -146
rect 264 -149 266 -146
rect 280 -149 282 -146
rect 296 -149 298 -146
rect 315 -149 317 -146
rect 331 -149 333 -146
rect 347 -149 349 -146
rect 363 -149 365 -146
rect 382 -149 384 -146
rect 398 -149 400 -146
rect 414 -149 416 -146
rect 430 -149 432 -146
rect 446 -149 448 -146
rect 462 -149 464 -146
rect 478 -149 480 -146
rect 494 -149 496 -146
rect 510 -149 512 -146
rect 528 -149 530 -146
rect 547 -149 549 -146
rect 567 -149 569 -146
rect 30 -194 32 -158
rect 46 -194 48 -158
rect 62 -194 64 -158
rect 83 -194 85 -158
rect 102 -194 104 -158
rect 122 -194 124 -158
rect 141 -194 143 -158
rect 232 -194 234 -158
rect 248 -194 250 -158
rect 264 -194 266 -158
rect 280 -194 282 -158
rect 296 -194 298 -158
rect 315 -194 317 -158
rect 331 -194 333 -158
rect 347 -194 349 -158
rect 363 -194 365 -158
rect 382 -194 384 -158
rect 398 -194 400 -158
rect 414 -194 416 -158
rect 430 -194 432 -158
rect 446 -194 448 -158
rect 462 -194 464 -158
rect 478 -194 480 -158
rect 494 -194 496 -158
rect 510 -194 512 -158
rect 528 -194 530 -158
rect 547 -194 549 -158
rect 567 -194 569 -158
rect 30 -201 32 -198
rect 46 -201 48 -198
rect 62 -201 64 -198
rect 83 -201 85 -198
rect 102 -201 104 -198
rect 122 -201 124 -198
rect 141 -201 143 -198
rect 232 -201 234 -198
rect 248 -201 250 -198
rect 264 -201 266 -198
rect 280 -201 282 -198
rect 296 -201 298 -198
rect 315 -201 317 -198
rect 331 -201 333 -198
rect 347 -201 349 -198
rect 363 -201 365 -198
rect 382 -201 384 -198
rect 398 -201 400 -198
rect 414 -201 416 -198
rect 430 -201 432 -198
rect 446 -201 448 -198
rect 462 -201 464 -198
rect 478 -201 480 -198
rect 494 -201 496 -198
rect 510 -201 512 -198
rect 528 -201 530 -198
rect 547 -201 549 -198
rect 567 -201 569 -198
rect 29 -220 31 -217
rect 45 -220 47 -217
rect 61 -220 63 -217
rect 82 -220 84 -217
rect 101 -220 103 -217
rect 121 -220 123 -217
rect 140 -220 142 -217
rect 232 -220 234 -217
rect 248 -220 250 -217
rect 264 -220 266 -217
rect 280 -220 282 -217
rect 296 -220 298 -217
rect 312 -220 314 -217
rect 328 -220 330 -217
rect 344 -220 346 -217
rect 360 -220 362 -217
rect 376 -220 378 -217
rect 392 -220 394 -217
rect 412 -220 414 -217
rect 428 -220 430 -217
rect 444 -220 446 -217
rect 460 -220 462 -217
rect 477 -220 479 -217
rect 493 -220 495 -217
rect 509 -220 511 -217
rect 525 -220 527 -217
rect 541 -220 543 -217
rect 557 -220 559 -217
rect 573 -220 575 -217
rect 589 -220 591 -217
rect 605 -220 607 -217
rect 29 -265 31 -229
rect 45 -265 47 -229
rect 61 -265 63 -229
rect 82 -265 84 -229
rect 101 -265 103 -229
rect 121 -265 123 -229
rect 140 -265 142 -229
rect 232 -265 234 -229
rect 248 -265 250 -229
rect 264 -265 266 -229
rect 280 -265 282 -229
rect 296 -265 298 -229
rect 312 -265 314 -229
rect 328 -265 330 -229
rect 344 -265 346 -229
rect 360 -265 362 -229
rect 376 -265 378 -229
rect 392 -265 394 -229
rect 412 -265 414 -229
rect 428 -265 430 -229
rect 444 -265 446 -229
rect 460 -265 462 -229
rect 477 -265 479 -229
rect 493 -265 495 -229
rect 509 -265 511 -229
rect 525 -265 527 -229
rect 541 -265 543 -229
rect 557 -265 559 -229
rect 573 -265 575 -229
rect 589 -265 591 -229
rect 605 -265 607 -229
rect 29 -272 31 -269
rect 45 -272 47 -269
rect 61 -272 63 -269
rect 82 -272 84 -269
rect 101 -272 103 -269
rect 121 -272 123 -269
rect 140 -272 142 -269
rect 232 -272 234 -269
rect 248 -272 250 -269
rect 264 -272 266 -269
rect 280 -272 282 -269
rect 296 -272 298 -269
rect 312 -272 314 -269
rect 328 -272 330 -269
rect 344 -272 346 -269
rect 360 -272 362 -269
rect 376 -272 378 -269
rect 392 -272 394 -269
rect 412 -272 414 -269
rect 428 -272 430 -269
rect 444 -272 446 -269
rect 460 -272 462 -269
rect 477 -272 479 -269
rect 493 -272 495 -269
rect 509 -272 511 -269
rect 525 -272 527 -269
rect 541 -272 543 -269
rect 557 -272 559 -269
rect 573 -272 575 -269
rect 589 -272 591 -269
rect 605 -272 607 -269
<< polycontact >>
rect 26 -29 30 -25
rect 42 -38 46 -34
rect 58 -29 62 -25
rect 79 -29 83 -25
rect 98 -38 102 -34
rect 118 -29 122 -25
rect 137 -48 141 -44
rect 219 -43 223 -38
rect 235 -35 239 -31
rect 251 -28 255 -24
rect 267 -29 271 -25
rect 287 -48 291 -44
rect 302 -39 307 -34
rect 318 -35 323 -30
rect 336 -28 341 -24
rect 356 -40 360 -35
rect 376 -49 380 -44
rect 26 -100 30 -96
rect 42 -109 46 -105
rect 58 -100 62 -96
rect 79 -100 83 -96
rect 98 -109 102 -105
rect 118 -100 122 -96
rect 137 -119 141 -115
rect 217 -101 221 -96
rect 237 -101 241 -96
rect 253 -120 257 -115
rect 269 -101 273 -97
rect 285 -105 289 -100
rect 301 -120 305 -115
rect 317 -101 321 -97
rect 336 -101 340 -96
rect 355 -119 359 -114
rect 371 -102 375 -97
rect 386 -110 391 -105
rect 402 -110 407 -105
rect 418 -106 423 -101
rect 436 -99 441 -95
rect 456 -111 460 -106
rect 476 -120 480 -115
rect 506 -116 511 -111
rect 524 -99 529 -95
rect 544 -111 548 -106
rect 564 -120 568 -115
rect 26 -171 30 -167
rect 42 -180 46 -176
rect 58 -171 62 -167
rect 79 -171 83 -167
rect 98 -180 102 -176
rect 118 -171 122 -167
rect 137 -190 141 -186
rect 228 -182 232 -177
rect 244 -173 248 -168
rect 260 -191 264 -186
rect 276 -173 280 -168
rect 292 -171 296 -167
rect 311 -182 315 -177
rect 327 -191 331 -186
rect 343 -182 347 -177
rect 359 -173 363 -169
rect 378 -191 382 -186
rect 394 -191 398 -186
rect 410 -173 414 -169
rect 425 -182 430 -177
rect 441 -182 446 -177
rect 458 -173 462 -168
rect 473 -182 478 -177
rect 490 -189 494 -185
rect 505 -177 510 -172
rect 523 -170 528 -166
rect 543 -182 547 -177
rect 563 -191 567 -186
rect 25 -242 29 -238
rect 41 -251 45 -247
rect 57 -242 61 -238
rect 78 -242 82 -238
rect 97 -251 101 -247
rect 117 -242 121 -238
rect 136 -261 140 -257
rect 228 -244 232 -239
rect 244 -244 248 -239
rect 260 -244 264 -239
rect 276 -244 280 -239
rect 292 -257 296 -253
rect 308 -241 312 -237
rect 323 -241 328 -237
rect 338 -248 344 -244
rect 356 -257 360 -253
rect 371 -248 376 -244
rect 388 -241 392 -237
rect 408 -243 412 -238
rect 424 -257 428 -253
rect 439 -244 444 -239
rect 456 -241 460 -237
rect 473 -257 477 -253
rect 489 -253 493 -248
rect 505 -241 509 -237
rect 521 -241 525 -237
rect 537 -252 541 -247
rect 553 -262 557 -257
rect 568 -244 573 -239
rect 584 -262 589 -257
rect 601 -241 605 -237
<< metal1 >>
rect 19 0 24 4
rect 29 0 352 4
rect 25 -7 29 0
rect 41 -7 45 0
rect 57 -7 61 0
rect 78 -7 82 0
rect 117 -7 121 0
rect 218 -7 222 0
rect 234 -7 238 0
rect 250 -7 254 0
rect 266 -7 270 0
rect 302 -7 306 0
rect 318 -7 322 0
rect 336 -7 340 0
rect 355 -4 394 -1
rect 355 -7 359 -4
rect 375 -7 379 -4
rect 90 -16 97 -7
rect 129 -16 136 -7
rect 278 -16 286 -7
rect 33 -25 37 -16
rect 49 -25 53 -16
rect 14 -29 20 -25
rect 33 -29 58 -25
rect 14 -38 36 -34
rect 49 -52 53 -29
rect 65 -43 69 -16
rect 105 -25 109 -16
rect 86 -29 118 -25
rect 65 -52 69 -49
rect 86 -52 90 -29
rect 105 -52 109 -29
rect 144 -31 148 -16
rect 226 -24 230 -16
rect 242 -24 246 -16
rect 226 -28 251 -24
rect 258 -25 262 -16
rect 144 -34 194 -31
rect 125 -35 194 -34
rect 125 -38 148 -35
rect 199 -35 235 -31
rect 125 -52 129 -38
rect 137 -44 141 -43
rect 137 -49 141 -48
rect 144 -52 148 -38
rect 208 -43 219 -38
rect 242 -52 246 -28
rect 258 -29 267 -25
rect 258 -52 262 -29
rect 294 -34 298 -16
rect 274 -39 302 -34
rect 310 -35 314 -16
rect 274 -52 278 -39
rect 294 -52 298 -39
rect 310 -40 318 -35
rect 310 -52 314 -40
rect 326 -44 330 -16
rect 344 -45 348 -16
rect 363 -19 367 -16
rect 363 -29 367 -24
rect 383 -20 387 -16
rect 363 -32 387 -29
rect 363 -39 371 -36
rect 363 -45 367 -39
rect 344 -49 367 -45
rect 326 -52 330 -49
rect 344 -52 348 -49
rect 363 -52 367 -49
rect 383 -52 387 -32
rect 37 -56 41 -52
rect 230 -56 234 -52
rect 25 -60 29 -56
rect 19 -64 36 -60
rect 57 -60 61 -56
rect 78 -60 82 -56
rect 97 -60 101 -56
rect 117 -60 121 -56
rect 136 -60 140 -56
rect 218 -60 222 -56
rect 250 -60 254 -56
rect 266 -60 270 -56
rect 286 -60 290 -56
rect 302 -60 306 -56
rect 318 -60 322 -56
rect 336 -60 340 -56
rect 355 -60 359 -56
rect 375 -60 379 -56
rect 391 -60 394 -4
rect 41 -64 350 -60
rect 355 -64 394 -60
rect 19 -71 24 -67
rect 29 -70 447 -67
rect 509 -70 540 -67
rect 29 -71 451 -70
rect 504 -71 540 -70
rect 25 -78 29 -72
rect 41 -78 45 -71
rect 57 -78 61 -71
rect 78 -78 82 -71
rect 117 -78 121 -71
rect 216 -78 220 -71
rect 236 -78 240 -71
rect 252 -78 256 -71
rect 268 -78 272 -71
rect 284 -78 288 -71
rect 300 -78 304 -71
rect 316 -78 320 -71
rect 335 -78 339 -71
rect 402 -78 406 -71
rect 418 -78 422 -71
rect 436 -78 440 -71
rect 455 -75 494 -72
rect 455 -78 459 -75
rect 475 -78 479 -75
rect 90 -87 97 -78
rect 129 -87 136 -78
rect 347 -87 354 -78
rect 366 -87 370 -78
rect 33 -96 37 -87
rect 49 -96 53 -87
rect 14 -100 20 -96
rect 33 -100 58 -96
rect 14 -109 36 -105
rect 49 -123 53 -100
rect 65 -114 69 -87
rect 105 -96 109 -87
rect 86 -100 118 -96
rect 65 -123 69 -120
rect 86 -123 90 -100
rect 105 -123 109 -100
rect 144 -102 148 -87
rect 125 -107 144 -105
rect 224 -106 228 -87
rect 244 -97 248 -87
rect 260 -97 264 -87
rect 276 -96 280 -87
rect 244 -101 269 -97
rect 292 -97 296 -87
rect 308 -97 312 -87
rect 244 -106 248 -101
rect 125 -109 148 -107
rect 125 -123 129 -109
rect 144 -123 148 -109
rect 224 -110 248 -106
rect 252 -120 253 -115
rect 260 -123 264 -101
rect 276 -123 280 -101
rect 292 -101 317 -97
rect 284 -106 289 -105
rect 308 -123 312 -101
rect 324 -114 328 -87
rect 378 -105 382 -87
rect 394 -105 398 -87
rect 343 -110 386 -105
rect 394 -110 402 -105
rect 410 -106 414 -87
rect 324 -123 328 -119
rect 343 -123 347 -110
rect 362 -123 366 -110
rect 378 -123 382 -110
rect 394 -123 398 -110
rect 410 -111 418 -106
rect 410 -123 414 -111
rect 426 -115 430 -87
rect 444 -116 448 -87
rect 463 -90 467 -87
rect 463 -100 467 -95
rect 483 -91 487 -87
rect 463 -103 487 -100
rect 463 -110 471 -107
rect 463 -116 467 -110
rect 444 -120 467 -116
rect 426 -123 430 -120
rect 444 -123 448 -120
rect 463 -123 467 -120
rect 483 -123 487 -103
rect 37 -127 41 -123
rect 228 -127 236 -123
rect 248 -127 252 -123
rect 296 -127 300 -123
rect 25 -131 29 -127
rect 19 -135 36 -131
rect 57 -131 61 -127
rect 78 -131 82 -127
rect 97 -131 101 -127
rect 117 -131 121 -127
rect 136 -131 140 -127
rect 216 -131 220 -127
rect 268 -131 272 -127
rect 284 -131 288 -127
rect 316 -131 320 -127
rect 335 -131 339 -127
rect 354 -131 358 -127
rect 370 -131 374 -127
rect 386 -131 390 -127
rect 402 -131 406 -127
rect 418 -131 422 -127
rect 436 -131 440 -127
rect 455 -131 459 -127
rect 475 -131 479 -127
rect 491 -131 494 -75
rect 506 -78 510 -71
rect 524 -78 528 -71
rect 543 -75 582 -72
rect 543 -78 547 -75
rect 563 -78 567 -75
rect 514 -115 518 -87
rect 532 -116 536 -87
rect 551 -90 555 -87
rect 551 -100 555 -95
rect 571 -91 575 -87
rect 551 -103 575 -100
rect 551 -110 559 -107
rect 551 -116 555 -110
rect 532 -120 555 -116
rect 514 -123 518 -120
rect 532 -123 536 -120
rect 551 -123 555 -120
rect 571 -123 575 -103
rect 506 -131 510 -127
rect 41 -135 450 -131
rect 455 -135 494 -131
rect 504 -135 513 -131
rect 524 -131 528 -127
rect 543 -131 547 -127
rect 563 -131 567 -127
rect 579 -131 582 -75
rect 518 -135 538 -131
rect 543 -135 582 -131
rect 19 -142 24 -138
rect 29 -142 539 -138
rect 25 -149 29 -143
rect 41 -149 45 -142
rect 57 -149 61 -142
rect 78 -149 82 -142
rect 117 -149 121 -142
rect 227 -149 231 -142
rect 243 -149 247 -142
rect 259 -149 263 -142
rect 275 -149 279 -142
rect 291 -149 295 -142
rect 310 -149 314 -142
rect 326 -149 330 -142
rect 342 -149 346 -142
rect 358 -149 362 -142
rect 377 -149 381 -142
rect 393 -149 397 -142
rect 409 -149 413 -142
rect 425 -149 429 -142
rect 489 -149 493 -142
rect 505 -149 509 -142
rect 523 -149 527 -142
rect 542 -146 581 -142
rect 542 -149 546 -146
rect 562 -149 566 -146
rect 90 -158 97 -149
rect 129 -158 136 -149
rect 437 -158 441 -149
rect 453 -158 457 -149
rect 469 -158 473 -149
rect 33 -167 37 -158
rect 49 -167 53 -158
rect 14 -171 20 -167
rect 33 -171 58 -167
rect 14 -180 36 -176
rect 49 -194 53 -171
rect 65 -185 69 -158
rect 105 -167 109 -158
rect 86 -171 118 -167
rect 65 -194 69 -191
rect 86 -194 90 -171
rect 105 -194 109 -171
rect 144 -172 148 -158
rect 235 -161 239 -158
rect 251 -161 255 -158
rect 267 -161 271 -158
rect 283 -161 287 -158
rect 235 -165 287 -161
rect 283 -167 287 -165
rect 125 -177 144 -176
rect 283 -171 292 -167
rect 299 -168 303 -158
rect 318 -161 322 -158
rect 334 -161 338 -158
rect 350 -161 354 -158
rect 318 -165 354 -161
rect 125 -180 148 -177
rect 125 -194 129 -180
rect 144 -194 148 -180
rect 283 -194 287 -171
rect 350 -169 354 -165
rect 350 -173 359 -169
rect 299 -194 303 -173
rect 350 -194 354 -173
rect 366 -177 370 -158
rect 385 -161 389 -158
rect 401 -161 405 -158
rect 385 -165 405 -161
rect 401 -169 405 -165
rect 401 -173 410 -169
rect 366 -194 370 -182
rect 401 -194 405 -173
rect 417 -177 421 -158
rect 417 -182 425 -177
rect 417 -194 421 -182
rect 481 -185 485 -158
rect 497 -177 501 -158
rect 497 -182 505 -177
rect 433 -189 490 -185
rect 433 -194 437 -189
rect 449 -194 453 -189
rect 465 -194 469 -189
rect 481 -194 485 -189
rect 497 -194 501 -182
rect 513 -186 517 -158
rect 531 -187 535 -158
rect 550 -161 554 -158
rect 550 -171 554 -166
rect 570 -162 574 -158
rect 550 -174 574 -171
rect 550 -181 558 -178
rect 550 -187 554 -181
rect 531 -191 554 -187
rect 513 -194 517 -191
rect 531 -194 535 -191
rect 550 -194 554 -191
rect 570 -194 574 -174
rect 37 -198 41 -194
rect 239 -198 243 -194
rect 255 -198 259 -194
rect 271 -198 275 -194
rect 322 -198 326 -194
rect 338 -198 342 -194
rect 389 -198 393 -194
rect 25 -202 29 -198
rect 19 -206 36 -202
rect 57 -202 61 -198
rect 78 -202 82 -198
rect 97 -202 101 -198
rect 117 -202 121 -198
rect 136 -202 140 -198
rect 227 -202 231 -198
rect 291 -202 295 -198
rect 310 -202 314 -198
rect 358 -202 362 -198
rect 377 -202 381 -198
rect 409 -202 413 -198
rect 425 -202 429 -198
rect 441 -202 445 -198
rect 457 -202 461 -198
rect 473 -202 477 -198
rect 489 -202 493 -198
rect 505 -202 509 -198
rect 41 -206 513 -202
rect 523 -202 527 -198
rect 542 -202 546 -198
rect 562 -202 566 -198
rect 578 -202 581 -146
rect 518 -206 537 -202
rect 542 -206 581 -202
rect 18 -213 24 -209
rect 29 -213 618 -209
rect 24 -220 28 -214
rect 40 -220 44 -213
rect 56 -220 60 -213
rect 77 -220 81 -213
rect 116 -220 120 -213
rect 227 -220 231 -213
rect 243 -220 247 -213
rect 259 -220 263 -213
rect 275 -220 279 -213
rect 291 -220 295 -213
rect 307 -220 311 -213
rect 323 -220 327 -213
rect 339 -220 343 -213
rect 355 -220 359 -213
rect 371 -220 375 -213
rect 407 -220 411 -213
rect 423 -220 427 -213
rect 439 -220 443 -213
rect 455 -220 459 -213
rect 472 -220 476 -213
rect 488 -220 492 -213
rect 504 -220 508 -213
rect 520 -220 524 -213
rect 600 -220 604 -213
rect 89 -229 96 -220
rect 128 -229 135 -220
rect 532 -229 536 -220
rect 548 -229 552 -220
rect 564 -229 568 -220
rect 580 -229 584 -220
rect 32 -238 36 -229
rect 48 -238 52 -229
rect 13 -242 19 -238
rect 32 -242 57 -238
rect 13 -251 35 -247
rect 48 -265 52 -242
rect 64 -256 68 -229
rect 104 -238 108 -229
rect 85 -242 117 -238
rect 64 -265 68 -262
rect 85 -265 89 -242
rect 104 -265 108 -242
rect 143 -247 147 -229
rect 235 -232 239 -229
rect 251 -232 255 -229
rect 267 -232 271 -229
rect 283 -232 287 -229
rect 299 -232 303 -229
rect 235 -236 303 -232
rect 299 -237 303 -236
rect 299 -241 308 -237
rect 124 -249 147 -247
rect 124 -251 296 -249
rect 124 -265 128 -251
rect 143 -253 296 -251
rect 143 -265 147 -253
rect 299 -265 303 -241
rect 315 -251 319 -229
rect 331 -232 335 -229
rect 347 -232 351 -229
rect 363 -232 367 -229
rect 379 -232 383 -229
rect 331 -236 383 -232
rect 379 -237 383 -236
rect 348 -251 353 -244
rect 379 -241 388 -237
rect 315 -254 353 -251
rect 315 -265 319 -254
rect 379 -265 383 -241
rect 395 -247 399 -229
rect 415 -232 419 -229
rect 431 -232 435 -229
rect 447 -232 451 -229
rect 415 -236 451 -232
rect 447 -237 451 -236
rect 463 -237 467 -229
rect 480 -232 484 -229
rect 496 -232 500 -229
rect 480 -236 500 -232
rect 496 -237 500 -236
rect 512 -237 516 -229
rect 592 -237 596 -229
rect 447 -241 456 -237
rect 417 -247 422 -244
rect 395 -250 422 -247
rect 395 -265 399 -250
rect 447 -265 451 -241
rect 463 -242 465 -237
rect 496 -241 505 -237
rect 512 -241 521 -237
rect 463 -265 467 -242
rect 496 -265 500 -241
rect 512 -265 516 -241
rect 592 -241 601 -237
rect 592 -265 596 -241
rect 608 -256 612 -229
rect 608 -260 616 -256
rect 608 -265 612 -260
rect 36 -269 40 -265
rect 239 -269 243 -265
rect 255 -269 259 -265
rect 271 -269 275 -265
rect 287 -269 291 -265
rect 335 -269 339 -265
rect 351 -269 355 -265
rect 367 -269 371 -265
rect 419 -269 423 -265
rect 435 -269 439 -265
rect 484 -269 488 -265
rect 24 -273 28 -269
rect 56 -273 60 -269
rect 77 -273 81 -269
rect 96 -273 100 -269
rect 116 -273 120 -269
rect 135 -273 139 -269
rect 227 -273 231 -269
rect 307 -273 311 -269
rect 323 -273 327 -269
rect 387 -273 391 -269
rect 407 -273 411 -269
rect 455 -273 459 -269
rect 472 -273 476 -269
rect 504 -273 508 -269
rect 520 -273 524 -269
rect 536 -273 540 -269
rect 552 -273 556 -269
rect 568 -273 572 -269
rect 584 -273 588 -269
rect 600 -273 604 -269
rect 18 -277 36 -273
rect 41 -277 615 -273
<< m2contact >>
rect 20 -30 26 -25
rect 36 -39 42 -34
rect 74 -30 79 -25
rect 65 -49 71 -43
rect 93 -39 98 -34
rect 194 -36 199 -31
rect 132 -49 137 -43
rect 203 -43 208 -38
rect 318 -40 323 -35
rect 336 -24 341 -19
rect 326 -49 331 -44
rect 362 -24 367 -19
rect 383 -25 388 -20
rect 351 -40 356 -35
rect 371 -40 376 -35
rect 371 -49 376 -44
rect 447 -70 452 -65
rect 504 -70 509 -65
rect 20 -101 26 -96
rect 36 -110 42 -105
rect 74 -101 79 -96
rect 93 -110 98 -105
rect 212 -101 217 -96
rect 144 -107 149 -102
rect 276 -101 281 -96
rect 331 -101 336 -96
rect 324 -119 329 -114
rect 350 -119 355 -114
rect 418 -111 423 -106
rect 436 -95 441 -90
rect 426 -120 431 -115
rect 462 -95 467 -90
rect 483 -96 488 -91
rect 451 -111 456 -106
rect 471 -111 476 -106
rect 471 -120 476 -115
rect 506 -111 511 -106
rect 524 -95 529 -90
rect 514 -120 519 -115
rect 550 -95 555 -90
rect 571 -96 576 -91
rect 539 -111 544 -106
rect 559 -111 564 -106
rect 559 -120 564 -115
rect 20 -172 26 -167
rect 36 -181 42 -176
rect 74 -172 79 -167
rect 93 -181 98 -176
rect 144 -177 149 -172
rect 271 -173 276 -168
rect 299 -173 304 -168
rect 366 -182 371 -177
rect 453 -173 458 -168
rect 436 -182 441 -177
rect 505 -182 510 -177
rect 523 -166 528 -161
rect 513 -191 518 -186
rect 549 -166 554 -161
rect 570 -167 575 -162
rect 538 -182 543 -177
rect 558 -182 563 -177
rect 558 -191 563 -186
rect 19 -243 25 -238
rect 35 -252 41 -247
rect 73 -243 78 -238
rect 92 -252 97 -247
rect 223 -244 228 -239
rect 239 -244 244 -239
rect 255 -244 260 -239
rect 271 -244 276 -239
rect 291 -262 296 -257
rect 338 -244 343 -239
rect 355 -262 360 -257
rect 434 -244 439 -239
rect 423 -262 428 -257
rect 465 -242 470 -237
rect 484 -253 489 -248
rect 472 -262 477 -257
rect 563 -244 568 -239
rect 579 -262 584 -257
<< metal2 >>
rect 341 -24 362 -19
rect 26 -30 74 -25
rect 371 -28 388 -25
rect 42 -39 93 -34
rect 371 -35 376 -28
rect 71 -49 132 -43
rect 137 -49 190 -43
rect 185 -51 190 -49
rect 26 -101 74 -96
rect 42 -110 93 -105
rect 149 -107 181 -102
rect 131 -120 132 -114
rect 137 -120 172 -114
rect 167 -124 172 -120
rect 167 -144 172 -129
rect 176 -115 181 -107
rect 26 -172 74 -167
rect 42 -181 93 -176
rect 149 -177 172 -172
rect 137 -191 163 -185
rect 167 -186 172 -177
rect 176 -177 181 -120
rect 185 -106 190 -56
rect 185 -153 190 -111
rect 194 -96 199 -36
rect 194 -168 199 -101
rect 323 -40 351 -37
rect 203 -74 208 -43
rect 331 -49 371 -44
rect 452 -70 504 -65
rect 203 -78 529 -74
rect 203 -96 208 -78
rect 231 -86 511 -82
rect 231 -96 237 -86
rect 441 -95 462 -90
rect 203 -101 212 -96
rect 281 -101 331 -96
rect 203 -160 208 -101
rect 471 -99 488 -96
rect 471 -106 476 -99
rect 423 -111 451 -108
rect 506 -106 511 -86
rect 524 -90 529 -78
rect 529 -95 550 -90
rect 559 -99 576 -96
rect 559 -106 564 -99
rect 511 -111 539 -108
rect 329 -119 350 -114
rect 431 -120 471 -115
rect 519 -120 559 -115
rect 203 -164 276 -160
rect 271 -168 276 -164
rect 528 -166 549 -161
rect 156 -195 161 -191
rect 25 -243 73 -238
rect 41 -252 92 -247
rect 156 -248 161 -200
rect 223 -229 228 -182
rect 223 -239 228 -234
rect 239 -239 244 -173
rect 304 -173 453 -168
rect 558 -170 575 -167
rect 255 -218 260 -191
rect 255 -239 260 -223
rect 271 -239 276 -173
rect 558 -177 563 -170
rect 371 -182 436 -177
rect 510 -182 538 -179
rect 338 -239 343 -182
rect 518 -191 558 -186
rect 389 -212 394 -191
rect 389 -217 439 -212
rect 434 -239 439 -217
rect 465 -229 568 -224
rect 465 -237 470 -229
rect 563 -239 568 -229
rect 156 -253 484 -248
rect 136 -257 147 -256
rect 136 -262 163 -257
rect 296 -262 335 -257
rect 340 -262 355 -257
rect 360 -262 423 -257
rect 428 -262 472 -257
rect 158 -267 163 -262
rect 579 -267 584 -262
rect 158 -272 584 -267
<< m3contact >>
rect 185 -56 190 -51
rect 167 -129 172 -124
rect 167 -149 172 -144
rect 176 -120 181 -115
rect 185 -111 190 -106
rect 185 -158 190 -153
rect 194 -101 199 -96
rect 194 -173 199 -168
rect 176 -182 181 -177
rect 167 -191 172 -186
rect 156 -200 161 -195
rect 223 -234 228 -229
rect 255 -223 260 -218
<< m123contact >>
rect 24 0 29 5
rect 336 -33 341 -28
rect 36 -64 41 -59
rect 24 -72 29 -67
rect 65 -120 71 -114
rect 132 -120 137 -114
rect 36 -135 41 -130
rect 24 -143 29 -138
rect 65 -191 71 -185
rect 132 -191 137 -185
rect 282 -49 287 -43
rect 231 -101 237 -96
rect 366 -102 371 -97
rect 436 -104 441 -99
rect 284 -111 289 -106
rect 247 -120 252 -115
rect 296 -120 301 -115
rect 513 -135 518 -130
rect 239 -173 244 -168
rect 223 -182 228 -177
rect 36 -206 41 -201
rect 24 -214 29 -209
rect 255 -191 260 -186
rect 523 -175 528 -170
rect 306 -182 311 -177
rect 338 -182 343 -177
rect 468 -182 473 -177
rect 322 -191 327 -186
rect 323 -237 328 -232
rect 373 -191 378 -186
rect 389 -191 394 -186
rect 513 -206 518 -201
rect 348 -244 353 -239
rect 371 -244 376 -239
rect 403 -243 408 -238
rect 417 -244 422 -239
rect 532 -252 537 -247
rect 64 -262 70 -256
rect 131 -262 136 -256
rect 548 -262 553 -257
rect 36 -278 41 -273
<< metal3 >>
rect 24 -67 29 0
rect 282 -51 287 -49
rect 190 -56 287 -51
rect 24 -138 29 -72
rect 24 -209 29 -143
rect 336 -64 341 -33
rect 36 -130 41 -64
rect 296 -68 341 -64
rect 199 -101 231 -96
rect 190 -111 284 -106
rect 71 -120 132 -114
rect 296 -115 301 -68
rect 181 -120 247 -115
rect 252 -120 296 -115
rect 366 -124 371 -102
rect 172 -129 371 -124
rect 436 -135 441 -104
rect 36 -201 41 -135
rect 361 -140 448 -135
rect 172 -149 394 -144
rect 190 -158 343 -153
rect 199 -173 239 -168
rect 338 -177 343 -158
rect 181 -182 223 -177
rect 228 -182 306 -177
rect 71 -191 132 -185
rect 389 -186 394 -149
rect 172 -191 255 -186
rect 260 -191 322 -186
rect 327 -191 356 -186
rect 361 -191 373 -186
rect 468 -195 473 -182
rect 161 -200 473 -195
rect 513 -201 518 -135
rect 523 -206 528 -175
rect 36 -273 41 -206
rect 260 -223 408 -218
rect 228 -232 328 -229
rect 228 -234 323 -232
rect 371 -239 376 -223
rect 403 -238 408 -223
rect 70 -262 131 -256
rect 348 -257 353 -244
rect 417 -247 422 -244
rect 417 -252 532 -247
rect 348 -262 548 -257
<< m234contact >>
rect 335 -262 340 -257
<< m4contact >>
rect 356 -140 361 -135
rect 356 -191 361 -186
rect 523 -211 528 -206
<< metal4 >>
rect 356 -186 361 -140
rect 335 -211 523 -206
rect 335 -257 340 -211
<< labels >>
rlabel metal1 613 -259 615 -257 7 c4
rlabel metal1 210 -42 212 -40 1 cr_in
rlabel metal1 502 -180 504 -178 1 c3
rlabel metal1 579 -183 581 -180 1 s3
rlabel metal1 391 -44 394 -41 1 s1
rlabel metal1 317 -40 320 -37 7 c1
rlabel metal1 29 -63 30 -62 1 gnd
rlabel metal1 80 2 91 3 5 vdd
rlabel metal3 112 -119 117 -116 1 g1
rlabel metal3 112 -190 117 -187 1 g2
rlabel metal3 111 -261 116 -258 1 g3
rlabel m2contact 144 -107 149 -102 1 p1
rlabel m2contact 144 -177 149 -172 1 p2
rlabel metal1 16 -29 19 -27 3 a0
rlabel metal1 17 -37 20 -35 3 b0
rlabel metal1 14 -100 17 -98 3 a1
rlabel metal1 15 -109 18 -107 3 b1
rlabel metal1 14 -171 17 -169 3 a2
rlabel metal1 15 -180 18 -178 3 b2
rlabel metal1 13 -242 16 -240 3 a3
rlabel metal1 13 -251 16 -249 3 b3
rlabel metal2 157 -48 160 -45 1 g0
rlabel metal1 158 -34 160 -32 1 p0
rlabel metal1 143 -249 147 -245 1 p3
rlabel metal1 417 -110 418 -109 1 c2
rlabel metal1 491 -114 494 -111 1 s2
rlabel metal1 579 -108 581 -106 1 s0
rlabel metal1 325 -107 327 -105 1 c2i2
rlabel metal1 277 -104 279 -102 1 c2i1
<< end >>
