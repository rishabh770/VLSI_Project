magic
tech scmos
timestamp 1638811332
<< error_p >>
rect 54 33 121 35
rect 54 31 60 33
rect 63 31 87 33
rect 90 31 120 33
rect 54 30 122 31
rect 54 28 55 30
rect 57 29 58 30
rect 59 29 61 30
rect 66 29 67 30
rect 68 29 73 30
rect 74 29 79 30
rect 56 28 61 29
rect 65 28 69 29
rect 72 28 73 29
rect 78 28 79 29
rect 54 26 61 28
rect 63 26 67 28
rect 71 27 73 28
rect 69 26 73 27
rect 56 25 61 26
rect 65 25 73 26
rect 77 26 79 28
rect 80 28 82 30
rect 84 29 85 30
rect 86 29 88 30
rect 92 29 100 30
rect 101 29 106 30
rect 107 29 112 30
rect 83 28 88 29
rect 80 26 88 28
rect 90 28 102 29
rect 105 28 106 29
rect 111 28 112 29
rect 90 27 94 28
rect 96 27 100 28
rect 104 27 106 28
rect 92 26 100 27
rect 102 26 106 27
rect 77 25 81 26
rect 83 25 88 26
rect 54 21 55 25
rect 57 22 58 25
rect 59 22 61 25
rect 66 22 67 25
rect 71 24 82 25
rect 72 22 73 24
rect 75 23 82 24
rect 77 22 82 23
rect 57 21 61 22
rect 54 19 61 21
rect 63 21 64 22
rect 66 21 68 22
rect 69 21 70 22
rect 72 21 74 22
rect 75 21 76 22
rect 78 21 82 22
rect 84 22 85 25
rect 86 22 88 25
rect 93 22 94 26
rect 98 25 106 26
rect 110 26 112 28
rect 113 28 115 30
rect 117 29 118 30
rect 119 29 121 30
rect 116 28 121 29
rect 113 26 121 28
rect 110 25 114 26
rect 116 25 121 26
rect 99 22 100 25
rect 104 24 115 25
rect 105 22 106 24
rect 108 23 115 24
rect 110 22 115 23
rect 84 21 88 22
rect 63 19 88 21
rect 90 21 91 22
rect 93 21 95 22
rect 96 21 97 22
rect 99 21 101 22
rect 102 21 103 22
rect 105 21 107 22
rect 108 21 109 22
rect 111 21 115 22
rect 117 22 118 25
rect 119 22 121 25
rect 117 21 121 22
rect 90 19 121 21
rect 54 18 122 19
rect 55 16 61 18
rect 62 16 81 18
rect 82 16 88 18
rect 89 16 114 18
rect 115 16 121 18
rect 56 15 57 16
rect 62 15 64 16
rect 65 15 66 16
rect 71 15 72 16
rect 77 15 78 16
rect 83 15 84 16
rect 89 15 91 16
rect 92 15 93 16
rect 98 15 99 16
rect 104 15 105 16
rect 110 15 111 16
rect 116 15 117 16
rect 57 4 60 6
rect 81 4 87 6
rect 139 4 151 6
rect 54 1 63 3
rect 54 0 55 1
rect 56 0 63 1
rect 65 1 104 3
rect 65 0 66 1
rect 67 0 104 1
rect 122 1 168 3
rect 122 0 123 1
rect 124 0 168 1
rect 56 -2 62 0
rect 67 -2 103 0
rect 123 -2 141 0
rect 143 -2 167 0
rect 54 -3 64 -2
rect 65 -3 105 -2
rect 123 -3 169 -2
rect 59 -4 60 -3
rect 61 -4 63 -3
rect 67 -4 83 -3
rect 84 -4 89 -3
rect 90 -4 95 -3
rect 58 -5 63 -4
rect 69 -5 85 -4
rect 88 -5 89 -4
rect 94 -5 95 -4
rect 55 -7 63 -5
rect 58 -8 63 -7
rect 59 -11 60 -8
rect 61 -11 63 -8
rect 70 -11 71 -5
rect 73 -6 77 -5
rect 79 -6 83 -5
rect 87 -6 89 -5
rect 75 -7 83 -6
rect 85 -7 89 -6
rect 76 -11 77 -7
rect 81 -8 89 -7
rect 93 -7 95 -5
rect 96 -5 98 -3
rect 100 -4 101 -3
rect 102 -4 104 -3
rect 123 -4 153 -3
rect 99 -5 104 -4
rect 125 -5 149 -4
rect 152 -5 153 -4
rect 154 -5 156 -3
rect 158 -4 159 -3
rect 160 -4 163 -3
rect 164 -4 165 -3
rect 166 -4 168 -3
rect 158 -5 168 -4
rect 96 -7 104 -5
rect 93 -8 97 -7
rect 99 -8 104 -7
rect 82 -11 83 -8
rect 87 -9 98 -8
rect 88 -11 89 -9
rect 91 -10 98 -9
rect 93 -11 98 -10
rect 56 -12 57 -11
rect 59 -12 63 -11
rect 56 -14 63 -12
rect 67 -12 68 -11
rect 70 -12 72 -11
rect 73 -12 74 -11
rect 76 -12 78 -11
rect 79 -12 80 -11
rect 82 -12 84 -11
rect 85 -12 86 -11
rect 88 -12 90 -11
rect 91 -12 92 -11
rect 94 -12 98 -11
rect 100 -11 101 -8
rect 102 -11 104 -8
rect 126 -11 127 -5
rect 128 -6 133 -5
rect 134 -6 168 -5
rect 130 -9 131 -8
rect 132 -9 133 -6
rect 138 -7 168 -6
rect 134 -9 136 -7
rect 130 -10 136 -9
rect 138 -10 139 -7
rect 140 -8 144 -7
rect 140 -10 142 -8
rect 146 -9 147 -7
rect 148 -8 150 -7
rect 148 -9 151 -8
rect 152 -9 153 -7
rect 154 -9 156 -7
rect 158 -9 159 -7
rect 160 -8 168 -7
rect 160 -9 162 -8
rect 146 -10 156 -9
rect 157 -10 162 -9
rect 164 -10 165 -8
rect 129 -11 165 -10
rect 166 -11 168 -8
rect 100 -12 104 -11
rect 67 -14 104 -12
rect 123 -12 124 -11
rect 126 -12 128 -11
rect 129 -12 168 -11
rect 123 -14 142 -12
rect 143 -14 168 -12
rect 54 -15 56 -14
rect 55 -17 56 -15
rect 57 -15 64 -14
rect 65 -15 67 -14
rect 57 -17 63 -15
rect 66 -17 67 -15
rect 68 -15 105 -14
rect 121 -15 123 -14
rect 124 -15 169 -14
rect 68 -17 97 -15
rect 98 -17 104 -15
rect 124 -17 135 -15
rect 136 -17 143 -15
rect 144 -17 149 -15
rect 150 -17 155 -15
rect 156 -17 161 -15
rect 162 -17 168 -15
rect 58 -18 59 -17
rect 69 -18 70 -17
rect 75 -18 76 -17
rect 81 -18 82 -17
rect 87 -18 88 -17
rect 93 -18 94 -17
rect 99 -18 100 -17
rect 125 -18 126 -17
rect 131 -18 132 -17
rect 137 -18 138 -17
rect 145 -18 146 -17
rect 151 -18 152 -17
rect 157 -18 158 -17
rect 163 -18 164 -17
rect 72 -26 78 -24
rect 96 -26 102 -24
rect 152 -26 158 -24
rect -13 -28 0 -26
rect -13 -29 -12 -28
rect -11 -31 0 -28
rect -13 -32 0 -31
rect 54 -29 59 -26
rect 60 -29 87 -26
rect 88 -29 109 -26
rect 140 -28 151 -26
rect 140 -29 141 -28
rect 142 -29 151 -28
rect 152 -29 169 -26
rect 54 -31 58 -29
rect 62 -31 86 -29
rect 90 -31 108 -29
rect 142 -31 165 -29
rect 166 -31 169 -29
rect 54 -32 110 -31
rect 140 -32 169 -31
rect -11 -33 -7 -32
rect -3 -33 -1 -32
rect 55 -33 56 -32
rect 57 -33 59 -32
rect 65 -33 66 -32
rect -9 -34 -1 -33
rect -8 -39 -7 -34
rect -5 -35 -1 -34
rect -3 -36 0 -35
rect -2 -39 -1 -36
rect 54 -37 59 -33
rect 64 -34 66 -33
rect 71 -34 72 -32
rect 77 -34 78 -32
rect 62 -36 66 -34
rect 70 -35 72 -34
rect 68 -36 72 -35
rect 64 -37 72 -36
rect 76 -36 78 -34
rect 79 -34 81 -32
rect 83 -33 84 -32
rect 85 -33 87 -32
rect 82 -34 87 -33
rect 93 -34 94 -32
rect 99 -34 100 -32
rect 79 -36 87 -34
rect 92 -35 94 -34
rect 76 -37 80 -36
rect 82 -37 87 -36
rect 90 -37 94 -35
rect 98 -36 100 -34
rect 101 -34 103 -32
rect 105 -33 106 -32
rect 107 -33 109 -32
rect 104 -34 109 -33
rect 143 -33 144 -32
rect 145 -33 161 -32
rect 163 -33 164 -32
rect 143 -34 164 -33
rect 101 -36 109 -34
rect 142 -35 156 -34
rect 157 -35 164 -34
rect 142 -36 164 -35
rect 165 -36 169 -32
rect 98 -37 102 -36
rect 104 -37 109 -36
rect 144 -37 169 -36
rect -11 -41 -10 -40
rect -9 -41 0 -39
rect 55 -40 56 -37
rect 57 -40 59 -37
rect 65 -39 66 -37
rect 70 -38 81 -37
rect 71 -39 72 -38
rect 74 -39 81 -38
rect 55 -41 59 -40
rect -11 -43 0 -41
rect -13 -44 -11 -43
rect -12 -46 -11 -44
rect -10 -44 0 -43
rect -10 -46 -5 -44
rect -4 -46 0 -44
rect 54 -43 59 -41
rect 62 -41 63 -40
rect 64 -41 81 -39
rect 83 -40 84 -37
rect 85 -40 87 -37
rect 92 -38 103 -37
rect 93 -39 94 -38
rect 96 -39 103 -38
rect 83 -41 87 -40
rect 62 -43 87 -41
rect 90 -41 91 -40
rect 92 -41 103 -39
rect 105 -40 106 -37
rect 107 -40 109 -37
rect 143 -39 169 -37
rect 105 -41 109 -40
rect 90 -43 109 -41
rect 142 -41 143 -40
rect 145 -41 169 -39
rect 142 -43 169 -41
rect 54 -44 62 -43
rect 54 -46 59 -44
rect -9 -47 -8 -46
rect -3 -47 -2 -46
rect 54 -47 55 -46
rect 61 -47 62 -44
rect 63 -44 90 -43
rect 63 -46 68 -44
rect 69 -46 74 -44
rect 75 -46 80 -44
rect 81 -46 87 -44
rect 64 -47 65 -46
rect 70 -47 71 -46
rect 76 -47 77 -46
rect 82 -47 83 -46
rect 89 -47 90 -44
rect 91 -44 110 -43
rect 140 -44 142 -43
rect 91 -46 96 -44
rect 97 -46 102 -44
rect 103 -46 109 -44
rect 141 -46 142 -44
rect 143 -44 169 -43
rect 143 -46 148 -44
rect 149 -45 152 -44
rect 149 -46 151 -45
rect 155 -46 160 -44
rect 161 -46 166 -44
rect 167 -46 169 -44
rect 92 -47 93 -46
rect 98 -47 99 -46
rect 104 -47 105 -46
rect 144 -47 145 -46
rect 150 -47 151 -46
rect 156 -47 157 -46
rect 162 -47 163 -46
<< ntransistor >>
rect 44 18 45 19
rect 50 18 51 19
rect 56 18 57 19
rect 65 18 66 19
rect 71 18 72 19
rect 77 18 78 19
rect 83 18 84 19
rect 92 18 93 19
rect 98 18 99 19
rect 104 18 105 19
rect 110 18 111 19
rect 116 18 117 19
rect 58 -15 59 -14
rect 69 -15 70 -14
rect 75 -15 76 -14
rect 81 -15 82 -14
rect 87 -15 88 -14
rect 93 -15 94 -14
rect 99 -15 100 -14
rect 125 -15 126 -14
rect 131 -15 132 -14
rect 137 -15 138 -14
rect 145 -15 146 -14
rect 151 -15 152 -14
rect 157 -15 158 -14
rect 163 -15 164 -14
rect -9 -44 -8 -43
rect -3 -44 -2 -43
rect 3 -44 4 -43
rect 9 -44 10 -43
rect 15 -44 16 -43
rect 21 -44 22 -43
rect 30 -44 31 -43
rect 36 -44 37 -43
rect 42 -44 43 -43
rect 48 -44 49 -43
rect 54 -44 55 -43
rect 64 -44 65 -43
rect 70 -44 71 -43
rect 76 -44 77 -43
rect 82 -44 83 -43
rect 92 -44 93 -43
rect 98 -44 99 -43
rect 104 -44 105 -43
rect 144 -44 145 -43
rect 150 -44 151 -43
rect 156 -44 157 -43
rect 162 -44 163 -43
<< ptransistor >>
rect 44 30 45 31
rect 50 30 51 31
rect 56 30 57 31
rect 65 30 66 31
rect 71 30 72 31
rect 77 30 78 31
rect 83 30 84 31
rect 92 30 93 31
rect 98 30 99 31
rect 104 30 105 31
rect 110 30 111 31
rect 116 30 117 31
rect 58 -3 59 -2
rect 69 -3 70 -2
rect 75 -3 76 -2
rect 81 -3 82 -2
rect 87 -3 88 -2
rect 93 -3 94 -2
rect 99 -3 100 -2
rect 125 -3 126 -2
rect 131 -3 132 -2
rect 137 -3 138 -2
rect 145 -3 146 -2
rect 151 -3 152 -2
rect 157 -3 158 -2
rect 163 -3 164 -2
rect -9 -32 -8 -31
rect -3 -32 -2 -31
rect 3 -32 4 -31
rect 9 -32 10 -31
rect 15 -32 16 -31
rect 21 -32 22 -31
rect 30 -32 31 -31
rect 36 -32 37 -31
rect 42 -32 43 -31
rect 48 -32 49 -31
rect 54 -32 55 -31
rect 64 -32 65 -31
rect 70 -32 71 -31
rect 76 -32 77 -31
rect 82 -32 83 -31
rect 92 -32 93 -31
rect 98 -32 99 -31
rect 104 -32 105 -31
rect 144 -32 145 -31
rect 150 -32 151 -31
rect 156 -32 157 -31
rect 162 -32 163 -31
<< ndiffusion >>
rect 43 18 44 19
rect 45 18 46 19
rect 47 18 48 19
rect 49 18 50 19
rect 51 18 52 19
rect 53 18 54 19
rect 55 18 56 19
rect 57 18 58 19
rect 59 18 60 19
rect 64 18 65 19
rect 66 18 67 19
rect 68 18 69 19
rect 70 18 71 19
rect 72 18 73 19
rect 74 18 75 19
rect 76 18 77 19
rect 78 18 79 19
rect 80 18 81 19
rect 82 18 83 19
rect 84 18 85 19
rect 86 18 87 19
rect 91 18 92 19
rect 93 18 94 19
rect 95 18 96 19
rect 97 18 98 19
rect 99 18 100 19
rect 101 18 102 19
rect 103 18 104 19
rect 105 18 106 19
rect 107 18 108 19
rect 109 18 110 19
rect 111 18 112 19
rect 113 18 114 19
rect 115 18 116 19
rect 117 18 118 19
rect 119 18 120 19
rect 57 -15 58 -14
rect 59 -15 60 -14
rect 68 -15 69 -14
rect 70 -15 71 -14
rect 72 -15 73 -14
rect 74 -15 75 -14
rect 76 -15 77 -14
rect 78 -15 79 -14
rect 80 -15 81 -14
rect 82 -15 83 -14
rect 84 -15 85 -14
rect 86 -15 87 -14
rect 88 -15 89 -14
rect 90 -15 91 -14
rect 92 -15 93 -14
rect 94 -15 95 -14
rect 96 -15 97 -14
rect 98 -15 99 -14
rect 100 -15 101 -14
rect 102 -15 103 -14
rect 124 -15 125 -14
rect 126 -15 127 -14
rect 128 -15 129 -14
rect 130 -15 131 -14
rect 132 -15 133 -14
rect 134 -15 135 -14
rect 136 -15 137 -14
rect 138 -15 139 -14
rect 140 -15 141 -14
rect 144 -15 145 -14
rect 146 -15 147 -14
rect 148 -15 149 -14
rect 150 -15 151 -14
rect 152 -15 153 -14
rect 154 -15 155 -14
rect 156 -15 157 -14
rect 158 -15 159 -14
rect 160 -15 161 -14
rect 162 -15 163 -14
rect 164 -15 165 -14
rect 166 -15 167 -14
rect -10 -44 -9 -43
rect -8 -44 -7 -43
rect -6 -44 -5 -43
rect -4 -44 -3 -43
rect -2 -44 -1 -43
rect 0 -44 1 -43
rect 2 -44 3 -43
rect 4 -44 5 -43
rect 6 -44 7 -43
rect 8 -44 9 -43
rect 10 -44 11 -43
rect 12 -44 13 -43
rect 14 -44 15 -43
rect 16 -44 17 -43
rect 18 -44 19 -43
rect 20 -44 21 -43
rect 22 -44 23 -43
rect 24 -44 25 -43
rect 29 -44 30 -43
rect 31 -44 32 -43
rect 33 -44 34 -43
rect 35 -44 36 -43
rect 37 -44 38 -43
rect 39 -44 40 -43
rect 41 -44 42 -43
rect 43 -44 44 -43
rect 45 -44 46 -43
rect 47 -44 48 -43
rect 49 -44 50 -43
rect 51 -44 52 -43
rect 53 -44 54 -43
rect 55 -44 56 -43
rect 57 -44 58 -43
rect 63 -44 64 -43
rect 65 -44 66 -43
rect 67 -44 68 -43
rect 69 -44 70 -43
rect 71 -44 72 -43
rect 73 -44 74 -43
rect 75 -44 76 -43
rect 77 -44 78 -43
rect 79 -44 80 -43
rect 81 -44 82 -43
rect 83 -44 84 -43
rect 85 -44 86 -43
rect 91 -44 92 -43
rect 93 -44 94 -43
rect 95 -44 96 -43
rect 97 -44 98 -43
rect 99 -44 100 -43
rect 101 -44 102 -43
rect 103 -44 104 -43
rect 105 -44 106 -43
rect 107 -44 108 -43
rect 143 -44 144 -43
rect 145 -44 146 -43
rect 147 -44 148 -43
rect 149 -44 150 -43
rect 151 -44 152 -43
rect 153 -44 154 -43
rect 155 -44 156 -43
rect 157 -44 158 -43
rect 159 -44 160 -43
rect 161 -44 162 -43
rect 163 -44 164 -43
<< pdiffusion >>
rect 42 30 43 31
rect 45 30 46 31
rect 47 30 48 31
rect 49 30 50 31
rect 51 30 52 31
rect 53 30 54 31
rect 55 30 56 31
rect 57 30 58 31
rect 59 30 60 31
rect 64 30 65 31
rect 66 30 67 31
rect 68 30 69 31
rect 70 30 71 31
rect 72 30 73 31
rect 74 30 75 31
rect 76 30 77 31
rect 78 30 79 31
rect 80 30 81 31
rect 82 30 83 31
rect 84 30 85 31
rect 86 30 87 31
rect 91 30 92 31
rect 93 30 94 31
rect 95 30 96 31
rect 97 30 98 31
rect 99 30 100 31
rect 101 30 102 31
rect 103 30 104 31
rect 105 30 106 31
rect 107 30 108 31
rect 109 30 110 31
rect 111 30 112 31
rect 113 30 114 31
rect 115 30 116 31
rect 117 30 118 31
rect 119 30 120 31
rect 57 -3 58 -2
rect 59 -3 60 -2
rect 61 -3 62 -2
rect 68 -3 69 -2
rect 70 -3 71 -2
rect 72 -3 73 -2
rect 74 -3 75 -2
rect 76 -3 77 -2
rect 78 -3 79 -2
rect 80 -3 81 -2
rect 82 -3 83 -2
rect 84 -3 85 -2
rect 86 -3 87 -2
rect 88 -3 89 -2
rect 90 -3 91 -2
rect 92 -3 93 -2
rect 94 -3 95 -2
rect 96 -3 97 -2
rect 98 -3 99 -2
rect 100 -3 101 -2
rect 102 -3 103 -2
rect 123 -3 124 -2
rect 126 -3 127 -2
rect 128 -3 129 -2
rect 130 -3 131 -2
rect 132 -3 133 -2
rect 134 -3 135 -2
rect 136 -3 137 -2
rect 138 -3 139 -2
rect 140 -3 141 -2
rect 144 -3 145 -2
rect 146 -3 147 -2
rect 148 -3 149 -2
rect 150 -3 151 -2
rect 152 -3 153 -2
rect 154 -3 155 -2
rect 156 -3 157 -2
rect 158 -3 159 -2
rect 160 -3 161 -2
rect 162 -3 163 -2
rect 164 -3 165 -2
rect 166 -3 167 -2
rect -10 -32 -9 -31
rect -8 -32 -7 -31
rect -6 -32 -5 -31
rect -4 -32 -3 -31
rect -2 -32 -1 -31
rect 0 -32 1 -31
rect 2 -32 3 -31
rect 4 -32 5 -31
rect 6 -32 7 -31
rect 8 -32 9 -31
rect 10 -32 11 -31
rect 12 -32 13 -31
rect 14 -32 15 -31
rect 16 -32 17 -31
rect 18 -32 19 -31
rect 20 -32 21 -31
rect 22 -32 23 -31
rect 24 -32 25 -31
rect 29 -32 30 -31
rect 31 -32 32 -31
rect 33 -32 34 -31
rect 35 -32 36 -31
rect 37 -32 38 -31
rect 39 -32 40 -31
rect 41 -32 42 -31
rect 43 -32 44 -31
rect 45 -32 46 -31
rect 47 -32 48 -31
rect 49 -32 50 -31
rect 51 -32 52 -31
rect 53 -32 54 -31
rect 55 -32 56 -31
rect 57 -32 58 -31
rect 63 -32 64 -31
rect 65 -32 66 -31
rect 67 -32 68 -31
rect 69 -32 70 -31
rect 71 -32 72 -31
rect 73 -32 74 -31
rect 75 -32 76 -31
rect 77 -32 78 -31
rect 79 -32 80 -31
rect 81 -32 82 -31
rect 83 -32 84 -31
rect 85 -32 86 -31
rect 91 -32 92 -31
rect 93 -32 94 -31
rect 95 -32 96 -31
rect 97 -32 98 -31
rect 99 -32 100 -31
rect 101 -32 102 -31
rect 103 -32 104 -31
rect 105 -32 106 -31
rect 107 -32 108 -31
rect 143 -32 144 -31
rect 145 -32 146 -31
rect 147 -32 148 -31
rect 149 -32 150 -31
rect 151 -32 152 -31
rect 153 -32 154 -31
rect 155 -32 156 -31
rect 157 -32 158 -31
rect 159 -32 160 -31
rect 161 -32 162 -31
rect 163 -32 164 -31
<< ndcontact >>
rect 42 18 43 19
rect 46 18 47 19
rect 48 18 49 19
rect 52 18 53 19
rect 54 18 55 19
rect 58 18 59 19
rect 63 18 64 19
rect 67 18 68 19
rect 69 18 70 19
rect 73 18 74 19
rect 75 18 76 19
rect 79 18 80 19
rect 81 18 82 19
rect 85 18 86 19
rect 90 18 91 19
rect 94 18 95 19
rect 96 18 97 19
rect 100 18 101 19
rect 102 18 103 19
rect 106 18 107 19
rect 108 18 109 19
rect 112 18 113 19
rect 114 18 115 19
rect 118 18 119 19
rect 56 -15 57 -14
rect 60 -15 61 -14
rect 67 -15 68 -14
rect 71 -15 72 -14
rect 73 -15 74 -14
rect 77 -15 78 -14
rect 79 -15 80 -14
rect 83 -15 84 -14
rect 85 -15 86 -14
rect 89 -15 90 -14
rect 91 -15 92 -14
rect 95 -15 96 -14
rect 97 -15 98 -14
rect 101 -15 102 -14
rect 123 -15 124 -14
rect 127 -15 128 -14
rect 129 -15 130 -14
rect 133 -15 134 -14
rect 135 -15 136 -14
rect 139 -15 140 -14
rect 143 -15 144 -14
rect 147 -15 148 -14
rect 149 -15 150 -14
rect 153 -15 154 -14
rect 155 -15 156 -14
rect 159 -15 160 -14
rect 161 -15 162 -14
rect 165 -15 166 -14
rect -11 -44 -10 -43
rect -7 -44 -6 -43
rect -5 -44 -4 -43
rect -1 -44 0 -43
rect 1 -44 2 -43
rect 5 -44 6 -43
rect 7 -44 8 -43
rect 11 -44 12 -43
rect 13 -44 14 -43
rect 17 -44 18 -43
rect 19 -44 20 -43
rect 23 -44 24 -43
rect 28 -44 29 -43
rect 32 -44 33 -43
rect 34 -44 35 -43
rect 38 -44 39 -43
rect 40 -44 41 -43
rect 44 -44 45 -43
rect 46 -44 47 -43
rect 50 -44 51 -43
rect 52 -44 53 -43
rect 56 -44 57 -43
rect 62 -44 63 -43
rect 66 -44 67 -43
rect 68 -44 69 -43
rect 72 -44 73 -43
rect 74 -44 75 -43
rect 78 -44 79 -43
rect 80 -44 81 -43
rect 84 -44 85 -43
rect 90 -44 91 -43
rect 94 -44 95 -43
rect 96 -44 97 -43
rect 100 -44 101 -43
rect 102 -44 103 -43
rect 106 -44 107 -43
rect 142 -44 143 -43
rect 146 -44 147 -43
rect 148 -44 149 -43
rect 152 -44 153 -43
rect 154 -44 155 -43
rect 158 -44 159 -43
rect 160 -44 161 -43
rect 164 -44 165 -43
<< pdcontact >>
rect 43 30 44 31
rect 46 30 47 31
rect 48 30 49 31
rect 52 30 53 31
rect 54 30 55 31
rect 58 30 59 31
rect 63 30 64 31
rect 67 30 68 31
rect 69 30 70 31
rect 73 30 74 31
rect 75 30 76 31
rect 79 30 80 31
rect 81 30 82 31
rect 85 30 86 31
rect 90 30 91 31
rect 94 30 95 31
rect 96 30 97 31
rect 100 30 101 31
rect 102 30 103 31
rect 106 30 107 31
rect 108 30 109 31
rect 112 30 113 31
rect 114 30 115 31
rect 118 30 119 31
rect 44 28 45 29
rect 50 25 51 26
rect 56 25 57 26
rect 65 25 66 26
rect 71 24 72 25
rect 77 22 78 23
rect 83 25 84 26
rect 92 26 93 27
rect 98 25 99 26
rect 104 24 105 25
rect 110 22 111 23
rect 116 25 117 26
rect 56 -3 57 -2
rect 60 -3 61 -2
rect 67 -3 68 -2
rect 71 -3 72 -2
rect 73 -3 74 -2
rect 77 -3 78 -2
rect 79 -3 80 -2
rect 83 -3 84 -2
rect 85 -3 86 -2
rect 89 -3 90 -2
rect 91 -3 92 -2
rect 95 -3 96 -2
rect 97 -3 98 -2
rect 101 -3 102 -2
rect 124 -3 125 -2
rect 127 -3 128 -2
rect 129 -3 130 -2
rect 133 -3 134 -2
rect 135 -3 136 -2
rect 139 -3 140 -2
rect 143 -3 144 -2
rect 147 -3 148 -2
rect 149 -3 150 -2
rect 153 -3 154 -2
rect 155 -3 156 -2
rect 159 -3 160 -2
rect 161 -3 162 -2
rect 165 -3 166 -2
rect 58 -8 59 -7
rect 69 -5 70 -4
rect 75 -7 76 -6
rect 81 -8 82 -7
rect 87 -9 88 -8
rect 93 -11 94 -10
rect 99 -8 100 -7
rect -11 -32 -10 -31
rect -7 -32 -6 -31
rect -5 -32 -4 -31
rect -1 -32 0 -31
rect 1 -32 2 -31
rect 5 -32 6 -31
rect 7 -32 8 -31
rect 11 -32 12 -31
rect 13 -32 14 -31
rect 17 -32 18 -31
rect 19 -32 20 -31
rect 23 -32 24 -31
rect 28 -32 29 -31
rect 32 -32 33 -31
rect 34 -32 35 -31
rect 38 -32 39 -31
rect 40 -32 41 -31
rect 44 -32 45 -31
rect 46 -32 47 -31
rect 50 -32 51 -31
rect 52 -32 53 -31
rect 56 -32 57 -31
rect 62 -32 63 -31
rect 66 -32 67 -31
rect 68 -32 69 -31
rect 72 -32 73 -31
rect 74 -32 75 -31
rect 78 -32 79 -31
rect 80 -32 81 -31
rect 84 -32 85 -31
rect 90 -32 91 -31
rect 94 -32 95 -31
rect 96 -32 97 -31
rect 100 -32 101 -31
rect 102 -32 103 -31
rect 106 -32 107 -31
rect 142 -32 143 -31
rect 146 -32 147 -31
rect 148 -32 149 -31
rect 152 -32 153 -31
rect 154 -32 155 -31
rect 158 -32 159 -31
rect 160 -32 161 -31
rect 164 -32 165 -31
rect -9 -34 -8 -33
rect -3 -36 -2 -35
rect 3 -37 4 -36
rect 9 -38 10 -37
rect 15 -40 16 -39
rect 21 -37 22 -36
rect 30 -36 31 -35
rect 36 -37 37 -36
rect 42 -38 43 -37
rect 48 -40 49 -39
rect 54 -37 55 -36
rect 64 -37 65 -36
rect 70 -38 71 -37
rect 76 -40 77 -39
rect 82 -37 83 -36
rect 92 -38 93 -37
rect 98 -40 99 -39
rect 104 -37 105 -36
<< polysilicon >>
rect 44 31 45 32
rect 50 31 51 32
rect 56 31 57 32
rect 65 31 66 32
rect 71 31 72 32
rect 77 31 78 32
rect 83 31 84 32
rect 92 31 93 32
rect 98 31 99 32
rect 104 31 105 32
rect 110 31 111 32
rect 116 31 117 32
rect 44 29 45 30
rect 44 19 45 28
rect 50 26 51 30
rect 50 19 51 25
rect 56 26 57 30
rect 56 19 57 25
rect 65 26 66 30
rect 65 19 66 25
rect 71 25 72 30
rect 71 19 72 24
rect 77 23 78 30
rect 77 19 78 22
rect 83 26 84 30
rect 83 19 84 25
rect 92 27 93 30
rect 92 19 93 26
rect 98 26 99 30
rect 98 19 99 25
rect 104 25 105 30
rect 104 19 105 24
rect 110 23 111 30
rect 110 19 111 22
rect 116 26 117 30
rect 116 19 117 25
rect 44 17 45 18
rect 50 17 51 18
rect 56 17 57 18
rect 65 17 66 18
rect 71 17 72 18
rect 77 17 78 18
rect 83 17 84 18
rect 92 17 93 18
rect 98 17 99 18
rect 104 17 105 18
rect 110 17 111 18
rect 116 17 117 18
rect 58 -2 59 -1
rect 69 -2 70 -1
rect 75 -2 76 -1
rect 81 -2 82 -1
rect 87 -2 88 -1
rect 93 -2 94 -1
rect 99 -2 100 -1
rect 125 -2 126 -1
rect 131 -2 132 -1
rect 137 -2 138 -1
rect 145 -2 146 -1
rect 151 -2 152 -1
rect 157 -2 158 -1
rect 163 -2 164 -1
rect 58 -7 59 -3
rect 58 -14 59 -8
rect 69 -4 70 -3
rect 69 -14 70 -5
rect 75 -6 76 -3
rect 75 -14 76 -7
rect 81 -7 82 -3
rect 81 -14 82 -8
rect 87 -8 88 -3
rect 87 -14 88 -9
rect 93 -10 94 -3
rect 93 -14 94 -11
rect 99 -7 100 -3
rect 99 -14 100 -8
rect 125 -4 126 -3
rect 125 -14 126 -5
rect 131 -12 132 -3
rect 131 -14 132 -13
rect 137 -6 138 -3
rect 137 -14 138 -7
rect 145 -4 146 -3
rect 145 -14 146 -5
rect 151 -12 152 -3
rect 151 -14 152 -13
rect 157 -12 158 -3
rect 157 -14 158 -13
rect 163 -7 164 -3
rect 163 -14 164 -8
rect 58 -16 59 -15
rect 69 -16 70 -15
rect 75 -16 76 -15
rect 81 -16 82 -15
rect 87 -16 88 -15
rect 93 -16 94 -15
rect 99 -16 100 -15
rect 125 -16 126 -15
rect 131 -16 132 -15
rect 137 -16 138 -15
rect 145 -16 146 -15
rect 151 -16 152 -15
rect 157 -16 158 -15
rect 163 -16 164 -15
rect -9 -31 -8 -30
rect -3 -31 -2 -30
rect 3 -31 4 -30
rect 9 -31 10 -30
rect 15 -31 16 -30
rect 21 -31 22 -30
rect 30 -31 31 -30
rect 36 -31 37 -30
rect 42 -31 43 -30
rect 48 -31 49 -30
rect 54 -31 55 -30
rect 64 -31 65 -30
rect 70 -31 71 -30
rect 76 -31 77 -30
rect 82 -31 83 -30
rect 92 -31 93 -30
rect 98 -31 99 -30
rect 104 -31 105 -30
rect 144 -31 145 -30
rect 150 -31 151 -30
rect 156 -31 157 -30
rect 162 -31 163 -30
rect -9 -33 -8 -32
rect -9 -43 -8 -34
rect -3 -35 -2 -32
rect -3 -43 -2 -36
rect 3 -36 4 -32
rect 3 -43 4 -37
rect 9 -37 10 -32
rect 9 -43 10 -38
rect 15 -39 16 -32
rect 15 -43 16 -40
rect 21 -36 22 -32
rect 21 -43 22 -37
rect 30 -35 31 -32
rect 30 -43 31 -36
rect 36 -36 37 -32
rect 36 -43 37 -37
rect 42 -37 43 -32
rect 42 -43 43 -38
rect 48 -39 49 -32
rect 48 -43 49 -40
rect 54 -36 55 -32
rect 54 -43 55 -37
rect 64 -36 65 -32
rect 64 -43 65 -37
rect 70 -37 71 -32
rect 70 -43 71 -38
rect 76 -39 77 -32
rect 76 -43 77 -40
rect 82 -36 83 -32
rect 82 -43 83 -37
rect 92 -37 93 -32
rect 92 -43 93 -38
rect 98 -39 99 -32
rect 98 -43 99 -40
rect 104 -36 105 -32
rect 104 -43 105 -37
rect 144 -36 145 -32
rect 144 -43 145 -37
rect 150 -35 151 -32
rect 150 -43 151 -36
rect 156 -38 157 -32
rect 156 -43 157 -39
rect 162 -41 163 -32
rect 162 -43 163 -42
rect -9 -45 -8 -44
rect -3 -45 -2 -44
rect 3 -45 4 -44
rect 9 -45 10 -44
rect 15 -45 16 -44
rect 21 -45 22 -44
rect 30 -45 31 -44
rect 36 -45 37 -44
rect 42 -45 43 -44
rect 48 -45 49 -44
rect 54 -45 55 -44
rect 64 -45 65 -44
rect 70 -45 71 -44
rect 76 -45 77 -44
rect 82 -45 83 -44
rect 92 -45 93 -44
rect 98 -45 99 -44
rect 104 -45 105 -44
rect 144 -45 145 -44
rect 150 -45 151 -44
rect 156 -45 157 -44
rect 162 -45 163 -44
<< polycontact >>
rect 125 -5 126 -4
rect 131 -13 132 -12
rect 137 -7 138 -6
rect 145 -5 146 -4
rect 151 -13 152 -12
rect 157 -13 158 -12
rect 163 -8 164 -7
rect 144 -37 145 -36
rect 150 -36 151 -35
rect 156 -39 157 -38
rect 162 -42 163 -41
<< metal1 >>
rect 42 33 61 34
rect 62 33 88 34
rect 89 33 121 34
rect 43 31 44 33
rect 48 31 49 33
rect 54 31 55 33
rect 63 31 64 33
rect 69 31 70 33
rect 75 31 76 33
rect 81 31 82 33
rect 90 31 91 33
rect 96 31 97 33
rect 102 31 103 33
rect 108 31 109 33
rect 114 31 115 33
rect 46 29 47 30
rect 52 29 53 30
rect 42 28 44 29
rect 46 28 53 29
rect 52 26 53 28
rect 58 26 59 30
rect 67 29 68 30
rect 73 29 74 30
rect 79 29 80 30
rect 67 28 80 29
rect 79 26 80 28
rect 85 26 86 30
rect 94 29 95 30
rect 100 29 101 30
rect 106 29 107 30
rect 112 29 113 30
rect 94 28 113 29
rect 90 26 92 27
rect 112 26 113 28
rect 118 26 119 30
rect 48 25 50 26
rect 52 25 56 26
rect 58 25 60 26
rect 63 25 65 26
rect 79 25 83 26
rect 85 25 87 26
rect 96 25 98 26
rect 112 25 116 26
rect 118 25 120 26
rect 52 19 53 25
rect 58 19 59 25
rect 69 24 71 25
rect 75 22 77 23
rect 79 19 80 25
rect 85 19 86 25
rect 102 24 104 25
rect 108 22 110 23
rect 112 19 113 25
rect 118 19 119 25
rect 47 18 48 19
rect 68 18 69 19
rect 74 18 75 19
rect 95 18 96 19
rect 101 18 102 19
rect 107 18 108 19
rect 42 16 43 18
rect 54 16 55 18
rect 63 16 64 18
rect 81 16 82 18
rect 90 16 91 18
rect 114 16 115 18
rect 42 15 61 16
rect 62 15 88 16
rect 89 15 121 16
rect 55 0 63 1
rect 66 0 104 1
rect 123 0 168 1
rect 56 -2 57 0
rect 67 -2 68 0
rect 73 -2 74 0
rect 79 -2 80 0
rect 85 -2 86 0
rect 91 -2 92 0
rect 97 -2 98 0
rect 124 -2 125 0
rect 129 -2 130 0
rect 135 -2 136 0
rect 143 -2 144 0
rect 155 -2 156 0
rect 161 -2 162 0
rect 148 -3 149 -2
rect 60 -7 61 -3
rect 71 -4 72 -3
rect 77 -4 78 -3
rect 83 -4 84 -3
rect 89 -4 90 -3
rect 95 -4 96 -3
rect 67 -5 69 -4
rect 71 -5 96 -4
rect 73 -7 75 -6
rect 95 -7 96 -5
rect 101 -7 102 -3
rect 123 -5 124 -4
rect 127 -6 128 -3
rect 133 -4 134 -3
rect 133 -6 134 -5
rect 127 -7 137 -6
rect 139 -7 140 -3
rect 153 -4 154 -3
rect 147 -5 154 -4
rect 55 -8 58 -7
rect 60 -8 62 -7
rect 79 -8 81 -7
rect 95 -8 99 -7
rect 101 -8 103 -7
rect 60 -14 61 -8
rect 85 -9 87 -8
rect 91 -11 93 -10
rect 95 -14 96 -8
rect 101 -14 102 -8
rect 129 -13 130 -12
rect 133 -14 134 -7
rect 139 -14 140 -8
rect 147 -14 148 -5
rect 153 -12 154 -5
rect 159 -12 160 -3
rect 165 -7 166 -3
rect 165 -8 167 -7
rect 165 -12 166 -8
rect 153 -13 157 -12
rect 159 -13 166 -12
rect 153 -14 154 -13
rect 159 -14 160 -13
rect 165 -14 166 -13
rect 72 -15 73 -14
rect 78 -15 79 -14
rect 84 -15 85 -14
rect 90 -15 91 -14
rect 128 -15 129 -14
rect 56 -17 57 -15
rect 67 -17 68 -15
rect 97 -17 98 -15
rect 123 -17 124 -15
rect 135 -17 136 -15
rect 143 -17 144 -15
rect 149 -17 150 -15
rect 155 -17 156 -15
rect 161 -17 162 -15
rect 55 -18 63 -17
rect 66 -18 104 -17
rect 123 -18 168 -17
rect -12 -29 26 -28
rect 27 -29 59 -28
rect 61 -29 87 -28
rect 89 -29 109 -28
rect 141 -29 149 -28
rect -11 -31 -10 -29
rect 19 -31 20 -29
rect 28 -31 29 -29
rect 52 -31 53 -29
rect 62 -31 63 -29
rect 80 -31 81 -29
rect 90 -31 91 -29
rect 102 -31 103 -29
rect 142 -31 143 -29
rect 148 -31 149 -29
rect 154 -29 167 -28
rect 154 -31 155 -29
rect 160 -31 161 -29
rect -6 -32 -5 -31
rect 0 -32 1 -31
rect 6 -32 7 -31
rect 12 -32 13 -31
rect 33 -32 34 -31
rect 39 -32 40 -31
rect 45 -32 46 -31
rect 67 -32 68 -31
rect 73 -32 74 -31
rect 95 -32 96 -31
rect -11 -34 -9 -33
rect -5 -36 -3 -35
rect 17 -36 18 -32
rect 23 -36 24 -32
rect 28 -36 30 -35
rect 50 -36 51 -32
rect 56 -36 57 -32
rect 78 -36 79 -32
rect 84 -36 85 -32
rect 100 -36 101 -32
rect 106 -36 107 -32
rect 1 -37 3 -36
rect 17 -37 21 -36
rect 23 -37 25 -36
rect 34 -37 36 -36
rect 50 -37 54 -36
rect 56 -37 58 -36
rect 62 -37 64 -36
rect 78 -37 82 -36
rect 84 -37 86 -36
rect 100 -37 104 -36
rect 106 -37 108 -36
rect 142 -37 143 -36
rect 7 -38 9 -37
rect 13 -40 15 -39
rect 17 -41 18 -37
rect -7 -42 18 -41
rect -7 -43 -6 -42
rect -1 -43 0 -42
rect 5 -43 6 -42
rect 11 -43 12 -42
rect 17 -43 18 -42
rect 23 -43 24 -37
rect 40 -38 42 -37
rect 46 -40 48 -39
rect 50 -41 51 -37
rect 32 -42 51 -41
rect 32 -43 33 -42
rect 38 -43 39 -42
rect 44 -43 45 -42
rect 50 -43 51 -42
rect 56 -43 57 -37
rect 68 -38 70 -37
rect 74 -40 76 -39
rect 78 -41 79 -37
rect 66 -42 79 -41
rect 66 -43 67 -42
rect 72 -43 73 -42
rect 78 -43 79 -42
rect 84 -43 85 -37
rect 90 -38 92 -37
rect 96 -40 98 -39
rect 100 -41 101 -37
rect 94 -42 101 -41
rect 94 -43 95 -42
rect 100 -43 101 -42
rect 106 -43 107 -37
rect 146 -41 147 -32
rect 148 -36 149 -35
rect 146 -43 147 -42
rect 152 -40 153 -32
rect 158 -33 159 -32
rect 158 -36 159 -34
rect 164 -38 165 -32
rect 158 -39 165 -38
rect 166 -36 167 -29
rect 166 -37 168 -36
rect 158 -40 159 -39
rect 152 -41 159 -40
rect 152 -43 153 -41
rect 158 -43 159 -41
rect 164 -43 165 -41
rect -11 -46 -10 -44
rect -5 -46 -4 -44
rect 1 -46 2 -44
rect 7 -46 8 -44
rect 13 -46 14 -44
rect 19 -46 20 -44
rect 28 -46 29 -44
rect 34 -46 35 -44
rect 40 -46 41 -44
rect 46 -46 47 -44
rect 52 -46 53 -44
rect 62 -46 63 -44
rect 68 -46 69 -44
rect 74 -46 75 -44
rect 80 -46 81 -44
rect 90 -46 91 -44
rect 96 -46 97 -44
rect 102 -46 103 -44
rect 142 -46 143 -44
rect 148 -46 149 -44
rect 154 -46 155 -44
rect 160 -46 161 -44
rect 166 -46 167 -37
rect -12 -47 26 -46
rect 27 -47 59 -46
rect 61 -47 87 -46
rect 89 -47 109 -46
rect 141 -47 150 -46
rect 154 -47 167 -46
<< m2contact >>
rect 124 -5 125 -4
rect 144 -5 145 -4
rect 130 -13 131 -12
rect 139 -8 140 -7
rect 162 -8 163 -7
rect 150 -13 151 -12
rect 143 -37 144 -36
rect 149 -36 150 -35
rect 146 -42 147 -41
rect 158 -34 159 -33
rect 158 -37 159 -36
rect 155 -39 156 -38
rect 164 -41 165 -40
rect 161 -42 162 -41
<< metal2 >>
rect 49 36 55 37
rect 72 36 78 37
rect 102 35 108 36
rect 57 3 60 4
rect 81 3 87 4
rect 139 3 151 4
rect 125 -5 144 -4
rect 140 -8 162 -7
rect 131 -13 150 -12
rect 3 -27 9 -26
rect 40 -27 46 -26
rect 72 -27 78 -26
rect 96 -27 102 -26
rect 152 -27 158 -26
rect 149 -34 158 -33
rect 149 -35 150 -34
rect 159 -37 161 -36
rect 143 -38 144 -37
rect 160 -38 161 -37
rect 143 -39 155 -38
rect 160 -39 165 -38
rect 164 -40 165 -39
rect 147 -42 161 -41
<< labels >>
rlabel metal1 24 -37 25 -36 1 Output
rlabel metal1 -11 -34 -10 -33 1 In5
rlabel metal1 -5 -36 -4 -35 1 In4
rlabel metal1 1 -37 2 -36 1 In3
rlabel metal1 7 -38 8 -37 1 In2
rlabel metal1 13 -40 14 -39 1 In1
rlabel metal2 3 -27 9 -26 1 5-input_OR
rlabel metal1 57 -37 58 -36 1 Output
rlabel metal1 28 -36 29 -35 1 In4
rlabel metal1 34 -37 35 -36 1 In3
rlabel metal1 40 -38 41 -37 1 In2
rlabel metal1 46 -40 47 -39 1 In1
rlabel metal2 40 -27 46 -26 1 4-input_OR
rlabel metal1 85 -37 86 -36 1 Output
rlabel metal1 62 -37 63 -36 1 In3
rlabel metal1 68 -38 69 -37 1 In2
rlabel metal1 74 -40 75 -39 1 In1
rlabel metal2 72 -27 78 -26 1 3-input_OR
rlabel metal1 107 -37 108 -36 1 Output
rlabel metal1 90 -38 91 -37 1 In2
rlabel metal1 96 -40 97 -39 1 In1
rlabel metal2 96 -27 102 -26 1 2-input_OR
rlabel metal1 123 -5 124 -4 3 In2
rlabel metal1 129 -13 130 -12 1 In1
rlabel metal1 166 -8 167 -7 1 Output
rlabel metal2 139 3 151 4 5 P_G_Block
rlabel metal1 75 22 76 23 1 In1
rlabel metal1 69 24 70 25 1 In2
rlabel metal1 63 25 64 26 1 In3
rlabel metal1 86 25 87 26 1 Output
rlabel metal2 72 36 78 37 5 3-input_AND
rlabel metal1 48 25 49 26 1 In1
rlabel metal1 59 25 60 26 1 Output
rlabel metal1 42 28 43 29 3 In2
rlabel metal2 49 36 55 37 5 2-input_AND
rlabel metal1 119 25 120 26 1 Output
rlabel metal1 90 26 91 27 1 In4
rlabel metal1 96 25 97 26 1 In3
rlabel metal1 102 24 103 25 1 In2
rlabel metal1 108 22 109 23 1 In1
rlabel metal2 102 35 108 36 1 4-input_AND
rlabel metal1 102 -8 103 -7 1 Output
rlabel metal1 67 -5 68 -4 1 In5
rlabel metal1 73 -7 74 -6 1 In4
rlabel metal1 79 -8 80 -7 1 In3
rlabel metal1 85 -9 86 -8 1 In2
rlabel metal1 91 -11 92 -10 1 In1
rlabel metal2 81 3 87 4 5 5-input_AND
rlabel metal1 61 -8 62 -7 1 Output
rlabel metal1 55 -8 57 -7 3 In
rlabel space 55 3 58 4 4 Inverter
rlabel metal1 142 -37 143 -36 1 In1
rlabel metal1 167 -37 168 -36 1 Output
rlabel metal1 148 -36 149 -35 1 In2
rlabel metal2 152 -27 158 -26 1 XOR_PTL
<< end >>
